magic
tech sky130A
magscale 1 2
timestamp 1745758139
<< nwell >>
rect 1066 2159 5834 9286
<< obsli1 >>
rect 1104 2159 5796 9265
<< obsm1 >>
rect 842 2128 5796 9296
<< obsm2 >>
rect 846 1391 5410 9625
<< metal3 >>
rect 0 9528 800 9648
rect 6100 9528 6900 9648
rect 0 6808 800 6928
rect 6100 6808 6900 6928
rect 0 4088 800 4208
rect 6100 4088 6900 4208
rect 0 1368 800 1488
rect 6100 1368 6900 1488
<< obsm3 >>
rect 880 9448 6020 9621
rect 798 7008 6100 9448
rect 880 6728 6020 7008
rect 798 4288 6100 6728
rect 880 4008 6020 4288
rect 798 1568 6100 4008
rect 880 1395 6020 1568
<< metal4 >>
rect 1944 2128 2264 9296
rect 2604 2128 2924 9296
<< labels >>
rlabel metal4 s 2604 2128 2924 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 9528 800 9648 6 a[0]
port 3 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 a[1]
port 4 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 a[2]
port 5 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 a[3]
port 6 nsew signal input
rlabel metal3 s 6100 9528 6900 9648 6 out[0]
port 7 nsew signal output
rlabel metal3 s 6100 6808 6900 6928 6 out[1]
port 8 nsew signal output
rlabel metal3 s 6100 4088 6900 4208 6 out[2]
port 9 nsew signal output
rlabel metal3 s 6100 1368 6900 1488 6 out[3]
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 6900 11424
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 101610
string GDS_FILE /openlane/designs/projectweek1/runs/RUN_2025.04.27_12.48.29/results/signoff/twos_complement.magic.gds
string GDS_START 52898
<< end >>

