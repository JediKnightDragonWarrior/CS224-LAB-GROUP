magic
tech sky130A
magscale 1 2
timestamp 1746356697
<< nwell >>
rect 1066 2159 10894 13638
<< obsli1 >>
rect 1104 2159 10856 13617
<< obsm1 >>
rect 842 2128 10934 13648
<< obsm2 >>
rect 846 575 10930 15337
<< metal3 >>
rect 0 15240 800 15360
rect 0 14424 800 14544
rect 11200 14424 12000 14544
rect 0 13608 800 13728
rect 0 12792 800 12912
rect 11200 12520 12000 12640
rect 0 11976 800 12096
rect 0 11160 800 11280
rect 11200 10616 12000 10736
rect 0 10344 800 10464
rect 0 9528 800 9648
rect 0 8712 800 8832
rect 11200 8712 12000 8832
rect 0 7896 800 8016
rect 0 7080 800 7200
rect 11200 6808 12000 6928
rect 0 6264 800 6384
rect 0 5448 800 5568
rect 11200 4904 12000 5024
rect 0 4632 800 4752
rect 0 3816 800 3936
rect 0 3000 800 3120
rect 11200 3000 12000 3120
rect 0 2184 800 2304
rect 0 1368 800 1488
rect 11200 1096 12000 1216
rect 0 552 800 672
<< obsm3 >>
rect 880 15160 11200 15333
rect 798 14624 11200 15160
rect 880 14344 11120 14624
rect 798 13808 11200 14344
rect 880 13528 11200 13808
rect 798 12992 11200 13528
rect 880 12720 11200 12992
rect 880 12712 11120 12720
rect 798 12440 11120 12712
rect 798 12176 11200 12440
rect 880 11896 11200 12176
rect 798 11360 11200 11896
rect 880 11080 11200 11360
rect 798 10816 11200 11080
rect 798 10544 11120 10816
rect 880 10536 11120 10544
rect 880 10264 11200 10536
rect 798 9728 11200 10264
rect 880 9448 11200 9728
rect 798 8912 11200 9448
rect 880 8632 11120 8912
rect 798 8096 11200 8632
rect 880 7816 11200 8096
rect 798 7280 11200 7816
rect 880 7008 11200 7280
rect 880 7000 11120 7008
rect 798 6728 11120 7000
rect 798 6464 11200 6728
rect 880 6184 11200 6464
rect 798 5648 11200 6184
rect 880 5368 11200 5648
rect 798 5104 11200 5368
rect 798 4832 11120 5104
rect 880 4824 11120 4832
rect 880 4552 11200 4824
rect 798 4016 11200 4552
rect 880 3736 11200 4016
rect 798 3200 11200 3736
rect 880 2920 11120 3200
rect 798 2384 11200 2920
rect 880 2104 11200 2384
rect 798 1568 11200 2104
rect 880 1296 11200 1568
rect 880 1288 11120 1296
rect 798 1016 11120 1288
rect 798 752 11200 1016
rect 880 579 11200 752
<< metal4 >>
rect 2163 2128 2483 13648
rect 2823 2128 3143 13648
rect 4601 2128 4921 13648
rect 5261 2128 5581 13648
rect 7039 2128 7359 13648
rect 7699 2128 8019 13648
rect 9477 2128 9797 13648
rect 10137 2128 10457 13648
<< metal5 >>
rect 1056 12672 10904 12992
rect 1056 12012 10904 12332
rect 1056 9816 10904 10136
rect 1056 9156 10904 9476
rect 1056 6960 10904 7280
rect 1056 6300 10904 6620
rect 1056 4104 10904 4424
rect 1056 3444 10904 3764
<< labels >>
rlabel metal3 s 0 6264 800 6384 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 A[2]
port 3 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 A[4]
port 5 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 A[5]
port 6 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 A[6]
port 7 nsew signal input
rlabel metal3 s 0 552 800 672 6 A[7]
port 8 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 B[0]
port 9 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 B[1]
port 10 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 B[2]
port 11 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 B[3]
port 12 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 B[4]
port 13 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 B[5]
port 14 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 B[6]
port 15 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 B[7]
port 16 nsew signal input
rlabel metal4 s 2823 2128 3143 13648 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 5261 2128 5581 13648 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 7699 2128 8019 13648 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 10137 2128 10457 13648 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 4104 10904 4424 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 6960 10904 7280 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 9816 10904 10136 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 12672 10904 12992 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 2163 2128 2483 13648 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 13648 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 13648 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 13648 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 3444 10904 3764 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 6300 10904 6620 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 9156 10904 9476 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 12012 10904 12332 6 VPWR
port 18 nsew power bidirectional
rlabel metal3 s 0 15240 800 15360 6 opcode[0]
port 19 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 opcode[1]
port 20 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 opcode[2]
port 21 nsew signal input
rlabel metal3 s 11200 14424 12000 14544 6 out[0]
port 22 nsew signal output
rlabel metal3 s 11200 12520 12000 12640 6 out[1]
port 23 nsew signal output
rlabel metal3 s 11200 10616 12000 10736 6 out[2]
port 24 nsew signal output
rlabel metal3 s 11200 8712 12000 8832 6 out[3]
port 25 nsew signal output
rlabel metal3 s 11200 6808 12000 6928 6 out[4]
port 26 nsew signal output
rlabel metal3 s 11200 4904 12000 5024 6 out[5]
port 27 nsew signal output
rlabel metal3 s 11200 3000 12000 3120 6 out[6]
port 28 nsew signal output
rlabel metal3 s 11200 1096 12000 1216 6 out[7]
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 12000 16000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 852798
string GDS_FILE /openlane/designs/projectweek2/runs/RUN_2025.05.04_11.04.10/results/signoff/lab2.magic.gds
string GDS_START 304114
<< end >>

