VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO twos_complement
  CLASS BLOCK ;
  FOREIGN twos_complement ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.500 BY 57.120 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 46.480 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END a[3]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 47.640 34.500 48.240 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 34.040 34.500 34.640 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 20.440 34.500 21.040 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 6.840 34.500 7.440 ;
    END
  END out[3]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 29.170 46.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 28.980 46.325 ;
      LAYER met1 ;
        RECT 4.210 10.640 28.980 46.480 ;
      LAYER met2 ;
        RECT 4.230 6.955 27.050 48.125 ;
      LAYER met3 ;
        RECT 4.400 47.240 30.100 48.105 ;
        RECT 3.990 35.040 30.500 47.240 ;
        RECT 4.400 33.640 30.100 35.040 ;
        RECT 3.990 21.440 30.500 33.640 ;
        RECT 4.400 20.040 30.100 21.440 ;
        RECT 3.990 7.840 30.500 20.040 ;
        RECT 4.400 6.975 30.100 7.840 ;
  END
END twos_complement
END LIBRARY

