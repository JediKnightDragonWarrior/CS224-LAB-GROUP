magic
tech sky130A
magscale 1 2
timestamp 1746356700
<< checkpaint >>
rect -3932 -3380 15932 19292
<< viali >>
rect 10425 13481 10459 13515
rect 1409 13345 1443 13379
rect 1685 13277 1719 13311
rect 2329 13277 2363 13311
rect 3065 13277 3099 13311
rect 3617 13277 3651 13311
rect 10241 13277 10275 13311
rect 2789 13209 2823 13243
rect 2973 13209 3007 13243
rect 2513 13141 2547 13175
rect 3249 13141 3283 13175
rect 3433 13141 3467 13175
rect 2237 12937 2271 12971
rect 3341 12937 3375 12971
rect 5365 12937 5399 12971
rect 1593 12801 1627 12835
rect 1685 12801 1719 12835
rect 2421 12801 2455 12835
rect 2697 12801 2731 12835
rect 2789 12801 2823 12835
rect 3157 12801 3191 12835
rect 3341 12801 3375 12835
rect 5273 12801 5307 12835
rect 5549 12801 5583 12835
rect 6377 12801 6411 12835
rect 7021 12801 7055 12835
rect 7205 12801 7239 12835
rect 10241 12801 10275 12835
rect 1961 12733 1995 12767
rect 6653 12733 6687 12767
rect 2421 12665 2455 12699
rect 5733 12665 5767 12699
rect 1501 12597 1535 12631
rect 2053 12597 2087 12631
rect 2973 12597 3007 12631
rect 6745 12597 6779 12631
rect 6929 12597 6963 12631
rect 7021 12597 7055 12631
rect 10425 12597 10459 12631
rect 6837 12393 6871 12427
rect 4261 12325 4295 12359
rect 6101 12325 6135 12359
rect 6653 12325 6687 12359
rect 3341 12257 3375 12291
rect 5089 12257 5123 12291
rect 2053 12189 2087 12223
rect 2145 12189 2179 12223
rect 2421 12189 2455 12223
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 3801 12189 3835 12223
rect 3893 12189 3927 12223
rect 4445 12189 4479 12223
rect 4808 12199 4842 12233
rect 4997 12189 5031 12223
rect 5273 12189 5307 12223
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 5641 12189 5675 12223
rect 6282 12189 6316 12223
rect 6745 12189 6779 12223
rect 7021 12189 7055 12223
rect 7113 12189 7147 12223
rect 7205 12189 7239 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 8125 12189 8159 12223
rect 8217 12189 8251 12223
rect 8493 12189 8527 12223
rect 4077 12121 4111 12155
rect 4905 12121 4939 12155
rect 5181 12121 5215 12155
rect 7323 12121 7357 12155
rect 7849 12121 7883 12155
rect 7941 12121 7975 12155
rect 8309 12121 8343 12155
rect 3801 12053 3835 12087
rect 5917 12053 5951 12087
rect 6285 12053 6319 12087
rect 7573 12053 7607 12087
rect 8401 12053 8435 12087
rect 2145 11849 2179 11883
rect 3081 11849 3115 11883
rect 3249 11849 3283 11883
rect 4997 11849 5031 11883
rect 5273 11849 5307 11883
rect 6561 11849 6595 11883
rect 8953 11849 8987 11883
rect 1961 11781 1995 11815
rect 2881 11781 2915 11815
rect 5089 11781 5123 11815
rect 7297 11781 7331 11815
rect 9229 11781 9263 11815
rect 1593 11713 1627 11747
rect 2237 11713 2271 11747
rect 2513 11713 2547 11747
rect 3341 11713 3375 11747
rect 3617 11713 3651 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 4813 11713 4847 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 5641 11713 5675 11747
rect 5917 11713 5951 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 7113 11713 7147 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 7481 11713 7515 11747
rect 7573 11713 7607 11747
rect 7757 11713 7791 11747
rect 8217 11713 8251 11747
rect 8861 11713 8895 11747
rect 9045 11713 9079 11747
rect 9321 11713 9355 11747
rect 2605 11645 2639 11679
rect 4721 11645 4755 11679
rect 5733 11645 5767 11679
rect 8309 11645 8343 11679
rect 4629 11577 4663 11611
rect 8585 11577 8619 11611
rect 8677 11577 8711 11611
rect 1961 11509 1995 11543
rect 3065 11509 3099 11543
rect 3433 11509 3467 11543
rect 3801 11509 3835 11543
rect 4537 11509 4571 11543
rect 7021 11509 7055 11543
rect 7941 11509 7975 11543
rect 9413 11509 9447 11543
rect 9781 11509 9815 11543
rect 2421 11305 2455 11339
rect 3341 11305 3375 11339
rect 3525 11305 3559 11339
rect 5181 11305 5215 11339
rect 5549 11305 5583 11339
rect 7297 11305 7331 11339
rect 8401 11305 8435 11339
rect 9689 11305 9723 11339
rect 9873 11305 9907 11339
rect 1593 11237 1627 11271
rect 2145 11237 2179 11271
rect 5089 11237 5123 11271
rect 8217 11237 8251 11271
rect 9597 11237 9631 11271
rect 10241 11237 10275 11271
rect 3985 11169 4019 11203
rect 5273 11169 5307 11203
rect 6285 11169 6319 11203
rect 8958 11169 8992 11203
rect 1409 11101 1443 11135
rect 1777 11101 1811 11135
rect 1961 11101 1995 11135
rect 3065 11101 3099 11135
rect 3433 11101 3467 11135
rect 4077 11101 4111 11135
rect 4445 11101 4479 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 4813 11101 4847 11135
rect 4905 11101 4939 11135
rect 5181 11101 5215 11135
rect 6469 11101 6503 11135
rect 9045 11101 9079 11135
rect 9416 11101 9450 11135
rect 2237 11033 2271 11067
rect 2437 11033 2471 11067
rect 3341 11033 3375 11067
rect 4353 11033 4387 11067
rect 6653 11033 6687 11067
rect 7113 11033 7147 11067
rect 7313 11033 7347 11067
rect 7941 11033 7975 11067
rect 9873 11033 9907 11067
rect 2605 10965 2639 10999
rect 3157 10965 3191 10999
rect 7481 10965 7515 10999
rect 9413 10965 9447 10999
rect 4813 10761 4847 10795
rect 10425 10761 10459 10795
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 4261 10625 4295 10659
rect 4997 10625 5031 10659
rect 5089 10625 5123 10659
rect 5181 10625 5215 10659
rect 5365 10625 5399 10659
rect 5457 10625 5491 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 6101 10625 6135 10659
rect 7849 10625 7883 10659
rect 8125 10625 8159 10659
rect 8217 10625 8251 10659
rect 10241 10625 10275 10659
rect 4353 10557 4387 10591
rect 5549 10557 5583 10591
rect 6009 10557 6043 10591
rect 8033 10557 8067 10591
rect 1593 10489 1627 10523
rect 4629 10489 4663 10523
rect 1869 10421 1903 10455
rect 4353 10421 4387 10455
rect 7849 10421 7883 10455
rect 4905 10217 4939 10251
rect 5641 10217 5675 10251
rect 9229 10149 9263 10183
rect 8953 10081 8987 10115
rect 2237 10013 2271 10047
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 3065 10013 3099 10047
rect 4721 10013 4755 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 1501 9945 1535 9979
rect 1685 9945 1719 9979
rect 2605 9945 2639 9979
rect 5641 9945 5675 9979
rect 2421 9877 2455 9911
rect 9413 9877 9447 9911
rect 3249 9673 3283 9707
rect 4169 9673 4203 9707
rect 6561 9605 6595 9639
rect 6745 9605 6779 9639
rect 1409 9537 1443 9571
rect 1501 9537 1535 9571
rect 1961 9537 1995 9571
rect 2605 9537 2639 9571
rect 3065 9537 3099 9571
rect 3801 9537 3835 9571
rect 6653 9537 6687 9571
rect 8769 9537 8803 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 9873 9537 9907 9571
rect 10057 9537 10091 9571
rect 1685 9469 1719 9503
rect 2053 9469 2087 9503
rect 2513 9469 2547 9503
rect 3893 9469 3927 9503
rect 8861 9469 8895 9503
rect 9413 9469 9447 9503
rect 9597 9469 9631 9503
rect 1593 9401 1627 9435
rect 2973 9401 3007 9435
rect 6377 9401 6411 9435
rect 9137 9401 9171 9435
rect 2237 9333 2271 9367
rect 6929 9333 6963 9367
rect 9229 9333 9263 9367
rect 9965 9333 9999 9367
rect 2697 9129 2731 9163
rect 2789 9129 2823 9163
rect 4077 9129 4111 9163
rect 4721 9129 4755 9163
rect 6469 9129 6503 9163
rect 7941 9129 7975 9163
rect 2881 9061 2915 9095
rect 6929 9061 6963 9095
rect 10425 9061 10459 9095
rect 5641 8993 5675 9027
rect 9413 8993 9447 9027
rect 10241 8993 10275 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 3157 8925 3191 8959
rect 3985 8925 4019 8959
rect 4537 8925 4571 8959
rect 5738 8925 5772 8959
rect 5917 8925 5951 8959
rect 6193 8925 6227 8959
rect 6285 8925 6319 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 9321 8925 9355 8959
rect 9965 8925 9999 8959
rect 10149 8925 10183 8959
rect 10517 8925 10551 8959
rect 5365 8857 5399 8891
rect 5549 8857 5583 8891
rect 5641 8857 5675 8891
rect 6101 8857 6135 8891
rect 6929 8857 6963 8891
rect 9781 8857 9815 8891
rect 2329 8789 2363 8823
rect 3341 8789 3375 8823
rect 4445 8789 4479 8823
rect 6653 8789 6687 8823
rect 7389 8789 7423 8823
rect 7481 8789 7515 8823
rect 8125 8789 8159 8823
rect 9689 8789 9723 8823
rect 10241 8789 10275 8823
rect 7297 8585 7331 8619
rect 7481 8585 7515 8619
rect 10425 8585 10459 8619
rect 6101 8517 6135 8551
rect 6469 8517 6503 8551
rect 6653 8517 6687 8551
rect 8369 8517 8403 8551
rect 8585 8517 8619 8551
rect 4261 8449 4295 8483
rect 4445 8449 4479 8483
rect 4537 8449 4571 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 6745 8449 6779 8483
rect 7356 8449 7390 8483
rect 7757 8449 7791 8483
rect 8953 8449 8987 8483
rect 9045 8449 9079 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 7849 8381 7883 8415
rect 5089 8313 5123 8347
rect 6469 8313 6503 8347
rect 8125 8313 8159 8347
rect 8217 8313 8251 8347
rect 9229 8313 9263 8347
rect 4353 8245 4387 8279
rect 4813 8245 4847 8279
rect 4997 8245 5031 8279
rect 8401 8245 8435 8279
rect 5457 8041 5491 8075
rect 6745 8041 6779 8075
rect 2053 7973 2087 8007
rect 2145 7973 2179 8007
rect 7849 7973 7883 8007
rect 4353 7905 4387 7939
rect 4445 7905 4479 7939
rect 4721 7905 4755 7939
rect 4813 7905 4847 7939
rect 4997 7905 5031 7939
rect 6653 7905 6687 7939
rect 7205 7905 7239 7939
rect 7297 7905 7331 7939
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 2697 7837 2731 7871
rect 2881 7837 2915 7871
rect 2973 7837 3007 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 4905 7837 4939 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5733 7837 5767 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 7113 7769 7147 7803
rect 8033 7769 8067 7803
rect 2421 7701 2455 7735
rect 2513 7701 2547 7735
rect 3985 7701 4019 7735
rect 5181 7701 5215 7735
rect 7757 7701 7791 7735
rect 2329 7497 2363 7531
rect 5273 7429 5307 7463
rect 1409 7361 1443 7395
rect 1961 7361 1995 7395
rect 2697 7361 2731 7395
rect 3893 7361 3927 7395
rect 4077 7361 4111 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 4629 7361 4663 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 4997 7361 5031 7395
rect 5089 7361 5123 7395
rect 10241 7361 10275 7395
rect 2053 7293 2087 7327
rect 2421 7293 2455 7327
rect 1593 7225 1627 7259
rect 3985 7225 4019 7259
rect 5273 7225 5307 7259
rect 2513 7157 2547 7191
rect 2881 7157 2915 7191
rect 4261 7157 4295 7191
rect 10425 7157 10459 7191
rect 5641 6953 5675 6987
rect 9781 6953 9815 6987
rect 1961 6885 1995 6919
rect 9873 6885 9907 6919
rect 3249 6817 3283 6851
rect 4353 6817 4387 6851
rect 4445 6817 4479 6851
rect 5733 6817 5767 6851
rect 6193 6817 6227 6851
rect 8217 6817 8251 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 2605 6749 2639 6783
rect 2697 6749 2731 6783
rect 2973 6749 3007 6783
rect 3065 6749 3099 6783
rect 3341 6749 3375 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 4721 6749 4755 6783
rect 4905 6749 4939 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 5457 6749 5491 6783
rect 5917 6749 5951 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 7297 6749 7331 6783
rect 7481 6749 7515 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9505 6749 9539 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 10149 6749 10183 6783
rect 1961 6681 1995 6715
rect 2329 6681 2363 6715
rect 2789 6681 2823 6715
rect 5273 6681 5307 6715
rect 5365 6681 5399 6715
rect 9873 6681 9907 6715
rect 1593 6613 1627 6647
rect 1777 6613 1811 6647
rect 2053 6613 2087 6647
rect 4629 6613 4663 6647
rect 4813 6613 4847 6647
rect 7389 6613 7423 6647
rect 8217 6613 8251 6647
rect 8953 6613 8987 6647
rect 10057 6613 10091 6647
rect 3617 6409 3651 6443
rect 5917 6409 5951 6443
rect 8233 6409 8267 6443
rect 8401 6409 8435 6443
rect 3249 6341 3283 6375
rect 3801 6341 3835 6375
rect 7205 6341 7239 6375
rect 8033 6341 8067 6375
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 5825 6273 5859 6307
rect 6101 6273 6135 6307
rect 6377 6273 6411 6307
rect 7113 6273 7147 6307
rect 7297 6273 7331 6307
rect 7573 6273 7607 6307
rect 8493 6273 8527 6307
rect 8585 6273 8619 6307
rect 9045 6273 9079 6307
rect 9689 6273 9723 6307
rect 7481 6205 7515 6239
rect 8769 6205 8803 6239
rect 9137 6205 9171 6239
rect 9413 6205 9447 6239
rect 9781 6205 9815 6239
rect 10057 6205 10091 6239
rect 6101 6137 6135 6171
rect 6561 6137 6595 6171
rect 7941 6137 7975 6171
rect 8217 6069 8251 6103
rect 8493 6069 8527 6103
rect 1593 5865 1627 5899
rect 7573 5865 7607 5899
rect 5917 5797 5951 5831
rect 7757 5797 7791 5831
rect 7849 5797 7883 5831
rect 9229 5797 9263 5831
rect 2145 5729 2179 5763
rect 8953 5729 8987 5763
rect 1409 5661 1443 5695
rect 2053 5661 2087 5695
rect 5733 5661 5767 5695
rect 7849 5661 7883 5695
rect 8125 5661 8159 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 8769 5661 8803 5695
rect 9505 5661 9539 5695
rect 9873 5661 9907 5695
rect 9965 5661 9999 5695
rect 7389 5593 7423 5627
rect 7589 5593 7623 5627
rect 2421 5525 2455 5559
rect 8033 5525 8067 5559
rect 8309 5525 8343 5559
rect 9413 5525 9447 5559
rect 9781 5525 9815 5559
rect 4169 5321 4203 5355
rect 5273 5321 5307 5355
rect 6561 5321 6595 5355
rect 9045 5321 9079 5355
rect 2329 5253 2363 5287
rect 4445 5253 4479 5287
rect 4645 5253 4679 5287
rect 5641 5253 5675 5287
rect 6377 5253 6411 5287
rect 1593 5185 1627 5219
rect 1685 5185 1719 5219
rect 1869 5185 1903 5219
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2513 5185 2547 5219
rect 2605 5185 2639 5219
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 4905 5185 4939 5219
rect 5825 5185 5859 5219
rect 5917 5185 5951 5219
rect 6045 5185 6079 5219
rect 6653 5185 6687 5219
rect 9413 5185 9447 5219
rect 10241 5185 10275 5219
rect 4997 5117 5031 5151
rect 9321 5117 9355 5151
rect 1869 5049 1903 5083
rect 1961 5049 1995 5083
rect 4353 5049 4387 5083
rect 4813 5049 4847 5083
rect 6377 5049 6411 5083
rect 3157 4981 3191 5015
rect 4629 4981 4663 5015
rect 5089 4981 5123 5015
rect 5641 4981 5675 5015
rect 10425 4981 10459 5015
rect 1593 4777 1627 4811
rect 3525 4777 3559 4811
rect 5089 4777 5123 4811
rect 4445 4641 4479 4675
rect 5365 4641 5399 4675
rect 1409 4573 1443 4607
rect 3433 4573 3467 4607
rect 3617 4573 3651 4607
rect 4537 4573 4571 4607
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 3801 4505 3835 4539
rect 3985 4505 4019 4539
rect 4169 4505 4203 4539
rect 4905 4437 4939 4471
rect 3801 4233 3835 4267
rect 2421 4165 2455 4199
rect 1409 4097 1443 4131
rect 1777 4097 1811 4131
rect 1869 4097 1903 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 2513 4097 2547 4131
rect 2697 4097 2731 4131
rect 2789 4097 2823 4131
rect 3065 4097 3099 4131
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 4261 4097 4295 4131
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 5273 4097 5307 4131
rect 5365 4097 5399 4131
rect 5549 4097 5583 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 7573 4097 7607 4131
rect 7849 4097 7883 4131
rect 8033 4097 8067 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 2881 4029 2915 4063
rect 5181 4029 5215 4063
rect 6561 4029 6595 4063
rect 2053 3961 2087 3995
rect 5089 3961 5123 3995
rect 1593 3893 1627 3927
rect 2145 3893 2179 3927
rect 3341 3893 3375 3927
rect 5733 3893 5767 3927
rect 7021 3893 7055 3927
rect 7849 3893 7883 3927
rect 8125 3893 8159 3927
rect 4445 3689 4479 3723
rect 4905 3689 4939 3723
rect 5733 3689 5767 3723
rect 4813 3621 4847 3655
rect 8953 3621 8987 3655
rect 1685 3553 1719 3587
rect 2145 3553 2179 3587
rect 4997 3553 5031 3587
rect 6285 3553 6319 3587
rect 6837 3553 6871 3587
rect 7021 3553 7055 3587
rect 7205 3553 7239 3587
rect 8217 3553 8251 3587
rect 2237 3485 2271 3519
rect 4353 3485 4387 3519
rect 4721 3485 4755 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 6377 3485 6411 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7573 3485 7607 3519
rect 7665 3485 7699 3519
rect 8125 3485 8159 3519
rect 9137 3485 9171 3519
rect 9326 3463 9360 3497
rect 10241 3485 10275 3519
rect 1501 3417 1535 3451
rect 5089 3417 5123 3451
rect 5549 3417 5583 3451
rect 8953 3417 8987 3451
rect 9229 3417 9263 3451
rect 2605 3349 2639 3383
rect 5749 3349 5783 3383
rect 5917 3349 5951 3383
rect 6009 3349 6043 3383
rect 7849 3349 7883 3383
rect 8493 3349 8527 3383
rect 10425 3349 10459 3383
rect 1961 3145 1995 3179
rect 4169 3145 4203 3179
rect 5549 3145 5583 3179
rect 7205 3145 7239 3179
rect 8223 3145 8257 3179
rect 1685 3077 1719 3111
rect 7481 3077 7515 3111
rect 8125 3077 8159 3111
rect 1501 3009 1535 3043
rect 1777 3009 1811 3043
rect 3249 3009 3283 3043
rect 3709 3009 3743 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 4537 3009 4571 3043
rect 5181 3009 5215 3043
rect 6653 3009 6687 3043
rect 6745 3009 6779 3043
rect 6837 3009 6871 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 8401 3009 8435 3043
rect 3157 2941 3191 2975
rect 3801 2941 3835 2975
rect 4629 2941 4663 2975
rect 4905 2941 4939 2975
rect 5273 2941 5307 2975
rect 6469 2941 6503 2975
rect 3617 2873 3651 2907
rect 5273 2805 5307 2839
rect 1685 2465 1719 2499
rect 1409 2397 1443 2431
rect 10241 2397 10275 2431
rect 10425 2261 10459 2295
<< metal1 >>
rect 1104 13626 10856 13648
rect 1104 13574 2169 13626
rect 2221 13574 2233 13626
rect 2285 13574 2297 13626
rect 2349 13574 2361 13626
rect 2413 13574 2425 13626
rect 2477 13574 4607 13626
rect 4659 13574 4671 13626
rect 4723 13574 4735 13626
rect 4787 13574 4799 13626
rect 4851 13574 4863 13626
rect 4915 13574 7045 13626
rect 7097 13574 7109 13626
rect 7161 13574 7173 13626
rect 7225 13574 7237 13626
rect 7289 13574 7301 13626
rect 7353 13574 9483 13626
rect 9535 13574 9547 13626
rect 9599 13574 9611 13626
rect 9663 13574 9675 13626
rect 9727 13574 9739 13626
rect 9791 13574 10856 13626
rect 1104 13552 10856 13574
rect 10410 13472 10416 13524
rect 10468 13472 10474 13524
rect 1394 13336 1400 13388
rect 1452 13336 1458 13388
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 2280 13280 2329 13308
rect 2280 13268 2286 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 3602 13268 3608 13320
rect 3660 13268 3666 13320
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 8628 13280 10241 13308
rect 8628 13268 8634 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 2774 13200 2780 13252
rect 2832 13200 2838 13252
rect 2961 13243 3019 13249
rect 2961 13209 2973 13243
rect 3007 13240 3019 13243
rect 3510 13240 3516 13252
rect 3007 13212 3516 13240
rect 3007 13209 3019 13212
rect 2961 13203 3019 13209
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 1452 13144 2513 13172
rect 1452 13132 1458 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 3234 13132 3240 13184
rect 3292 13132 3298 13184
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 3384 13144 3433 13172
rect 3384 13132 3390 13144
rect 3421 13141 3433 13144
rect 3467 13141 3479 13175
rect 3421 13135 3479 13141
rect 1104 13082 10856 13104
rect 1104 13030 2829 13082
rect 2881 13030 2893 13082
rect 2945 13030 2957 13082
rect 3009 13030 3021 13082
rect 3073 13030 3085 13082
rect 3137 13030 5267 13082
rect 5319 13030 5331 13082
rect 5383 13030 5395 13082
rect 5447 13030 5459 13082
rect 5511 13030 5523 13082
rect 5575 13030 7705 13082
rect 7757 13030 7769 13082
rect 7821 13030 7833 13082
rect 7885 13030 7897 13082
rect 7949 13030 7961 13082
rect 8013 13030 10143 13082
rect 10195 13030 10207 13082
rect 10259 13030 10271 13082
rect 10323 13030 10335 13082
rect 10387 13030 10399 13082
rect 10451 13030 10856 13082
rect 1104 13008 10856 13030
rect 2222 12928 2228 12980
rect 2280 12928 2286 12980
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2648 12940 3341 12968
rect 2648 12928 2654 12940
rect 3329 12937 3341 12940
rect 3375 12937 3387 12971
rect 3329 12931 3387 12937
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 5353 12971 5411 12977
rect 5353 12968 5365 12971
rect 5040 12940 5365 12968
rect 5040 12928 5046 12940
rect 5353 12937 5365 12940
rect 5399 12937 5411 12971
rect 5353 12931 5411 12937
rect 3234 12900 3240 12912
rect 1596 12872 3240 12900
rect 1596 12841 1624 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1670 12792 1676 12844
rect 1728 12792 1734 12844
rect 1946 12724 1952 12776
rect 2004 12724 2010 12776
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2240 12628 2268 12872
rect 2406 12792 2412 12844
rect 2464 12792 2470 12844
rect 2700 12841 2728 12872
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 5276 12872 6316 12900
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2498 12724 2504 12776
rect 2556 12764 2562 12776
rect 2792 12764 2820 12795
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2924 12804 3157 12832
rect 2924 12792 2930 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 5276 12841 5304 12872
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 2556 12736 2820 12764
rect 2556 12724 2562 12736
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5552 12764 5580 12795
rect 6288 12776 6316 12872
rect 6362 12792 6368 12844
rect 6420 12792 6426 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 7926 12832 7932 12844
rect 7239 12804 7932 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 5224 12736 5580 12764
rect 5224 12724 5230 12736
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6328 12736 6653 12764
rect 6328 12724 6334 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 7024 12764 7052 12795
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 7374 12764 7380 12776
rect 7024 12736 7380 12764
rect 6641 12727 6699 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 5534 12696 5540 12708
rect 2455 12668 5540 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 8570 12696 8576 12708
rect 5767 12668 8576 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 8570 12656 8576 12668
rect 8628 12656 8634 12708
rect 2096 12600 2268 12628
rect 2961 12631 3019 12637
rect 2096 12588 2102 12600
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 4522 12628 4528 12640
rect 3007 12600 4528 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 6733 12631 6791 12637
rect 6733 12597 6745 12631
rect 6779 12628 6791 12631
rect 6822 12628 6828 12640
rect 6779 12600 6828 12628
rect 6779 12597 6791 12600
rect 6733 12591 6791 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7466 12628 7472 12640
rect 7055 12600 7472 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 10410 12588 10416 12640
rect 10468 12588 10474 12640
rect 1104 12538 10856 12560
rect 1104 12486 2169 12538
rect 2221 12486 2233 12538
rect 2285 12486 2297 12538
rect 2349 12486 2361 12538
rect 2413 12486 2425 12538
rect 2477 12486 4607 12538
rect 4659 12486 4671 12538
rect 4723 12486 4735 12538
rect 4787 12486 4799 12538
rect 4851 12486 4863 12538
rect 4915 12486 7045 12538
rect 7097 12486 7109 12538
rect 7161 12486 7173 12538
rect 7225 12486 7237 12538
rect 7289 12486 7301 12538
rect 7353 12486 9483 12538
rect 9535 12486 9547 12538
rect 9599 12486 9611 12538
rect 9663 12486 9675 12538
rect 9727 12486 9739 12538
rect 9791 12486 10856 12538
rect 1104 12464 10856 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 3326 12424 3332 12436
rect 2004 12396 3332 12424
rect 2004 12384 2010 12396
rect 1670 12316 1676 12368
rect 1728 12356 1734 12368
rect 2682 12356 2688 12368
rect 1728 12328 2688 12356
rect 1728 12316 1734 12328
rect 2038 12180 2044 12232
rect 2096 12180 2102 12232
rect 2148 12229 2176 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 2682 12220 2688 12232
rect 2464 12192 2688 12220
rect 2464 12180 2470 12192
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2884 12229 2912 12396
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4632 12396 6224 12424
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 4249 12359 4307 12365
rect 4249 12356 4261 12359
rect 4028 12328 4261 12356
rect 4028 12316 4034 12328
rect 4249 12325 4261 12328
rect 4295 12356 4307 12359
rect 4430 12356 4436 12368
rect 4295 12328 4436 12356
rect 4295 12325 4307 12328
rect 4249 12319 4307 12325
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 3326 12248 3332 12300
rect 3384 12248 3390 12300
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 3568 12260 4200 12288
rect 3568 12248 3574 12260
rect 4172 12232 4200 12260
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 1486 12112 1492 12164
rect 1544 12152 1550 12164
rect 1946 12152 1952 12164
rect 1544 12124 1952 12152
rect 1544 12112 1550 12124
rect 1946 12112 1952 12124
rect 2004 12152 2010 12164
rect 3068 12152 3096 12183
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3789 12223 3847 12229
rect 3789 12220 3801 12223
rect 3476 12192 3801 12220
rect 3476 12180 3482 12192
rect 3789 12189 3801 12192
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3878 12180 3884 12232
rect 3936 12180 3942 12232
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4212 12192 4445 12220
rect 4212 12180 4218 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 2004 12124 3096 12152
rect 2004 12112 2010 12124
rect 3602 12112 3608 12164
rect 3660 12152 3666 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3660 12124 4077 12152
rect 3660 12112 3666 12124
rect 4065 12121 4077 12124
rect 4111 12152 4123 12155
rect 4632 12152 4660 12396
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5902 12356 5908 12368
rect 4764 12328 5908 12356
rect 4764 12316 4770 12328
rect 4816 12239 4844 12328
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 4948 12260 5028 12288
rect 4948 12248 4954 12260
rect 4796 12233 4854 12239
rect 4796 12199 4808 12233
rect 4842 12199 4854 12233
rect 5000 12229 5028 12260
rect 5074 12248 5080 12300
rect 5132 12248 5138 12300
rect 5276 12229 5304 12328
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 6086 12316 6092 12368
rect 6144 12316 6150 12368
rect 5810 12288 5816 12300
rect 5368 12260 5816 12288
rect 4796 12193 4854 12199
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12189 5043 12223
rect 4985 12183 5043 12189
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 4111 12124 4660 12152
rect 4893 12155 4951 12161
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 4893 12121 4905 12155
rect 4939 12121 4951 12155
rect 4893 12115 4951 12121
rect 5169 12155 5227 12161
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 5368 12152 5396 12260
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5215 12124 5396 12152
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 4154 12084 4160 12096
rect 3835 12056 4160 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 4908 12084 4936 12115
rect 5460 12084 5488 12183
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5626 12180 5632 12232
rect 5684 12180 5690 12232
rect 6196 12220 6224 12396
rect 6822 12384 6828 12436
rect 6880 12384 6886 12436
rect 6641 12359 6699 12365
rect 6641 12325 6653 12359
rect 6687 12356 6699 12359
rect 6914 12356 6920 12368
rect 6687 12328 6920 12356
rect 6687 12325 6699 12328
rect 6641 12319 6699 12325
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 7742 12356 7748 12368
rect 7064 12328 7748 12356
rect 7064 12316 7070 12328
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 7984 12328 8524 12356
rect 7984 12316 7990 12328
rect 7208 12260 8432 12288
rect 6270 12223 6328 12229
rect 6270 12220 6282 12223
rect 6196 12192 6282 12220
rect 6270 12189 6282 12192
rect 6316 12220 6328 12223
rect 6316 12192 6408 12220
rect 6316 12189 6328 12192
rect 6270 12183 6328 12189
rect 6380 12152 6408 12192
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6604 12192 6745 12220
rect 6604 12180 6610 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7024 12152 7052 12183
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 7208 12229 7236 12260
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7558 12220 7564 12232
rect 7515 12192 7564 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 8168 12192 8217 12220
rect 8168 12180 8174 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 6380 12124 6960 12152
rect 7024 12124 7236 12152
rect 6932 12096 6960 12124
rect 4856 12056 5488 12084
rect 4856 12044 4862 12056
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 5684 12056 5917 12084
rect 5684 12044 5690 12056
rect 5905 12053 5917 12056
rect 5951 12053 5963 12087
rect 5905 12047 5963 12053
rect 6270 12044 6276 12096
rect 6328 12044 6334 12096
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 7208 12084 7236 12124
rect 7282 12112 7288 12164
rect 7340 12161 7346 12164
rect 7340 12155 7369 12161
rect 7357 12121 7369 12155
rect 7340 12115 7369 12121
rect 7837 12155 7895 12161
rect 7837 12121 7849 12155
rect 7883 12121 7895 12155
rect 7837 12115 7895 12121
rect 7340 12112 7346 12115
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7208 12056 7573 12084
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7852 12084 7880 12115
rect 7926 12112 7932 12164
rect 7984 12112 7990 12164
rect 8297 12155 8355 12161
rect 8297 12121 8309 12155
rect 8343 12121 8355 12155
rect 8297 12115 8355 12121
rect 8202 12084 8208 12096
rect 7852 12056 8208 12084
rect 7561 12047 7619 12053
rect 8202 12044 8208 12056
rect 8260 12084 8266 12096
rect 8312 12084 8340 12115
rect 8404 12093 8432 12260
rect 8496 12229 8524 12328
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8260 12056 8340 12084
rect 8389 12087 8447 12093
rect 8260 12044 8266 12056
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 9306 12084 9312 12096
rect 8435 12056 9312 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 1104 11994 10856 12016
rect 1104 11942 2829 11994
rect 2881 11942 2893 11994
rect 2945 11942 2957 11994
rect 3009 11942 3021 11994
rect 3073 11942 3085 11994
rect 3137 11942 5267 11994
rect 5319 11942 5331 11994
rect 5383 11942 5395 11994
rect 5447 11942 5459 11994
rect 5511 11942 5523 11994
rect 5575 11942 7705 11994
rect 7757 11942 7769 11994
rect 7821 11942 7833 11994
rect 7885 11942 7897 11994
rect 7949 11942 7961 11994
rect 8013 11942 10143 11994
rect 10195 11942 10207 11994
rect 10259 11942 10271 11994
rect 10323 11942 10335 11994
rect 10387 11942 10399 11994
rect 10451 11942 10856 11994
rect 1104 11920 10856 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 2498 11880 2504 11892
rect 2179 11852 2504 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 3069 11883 3127 11889
rect 3069 11880 3081 11883
rect 2740 11852 3081 11880
rect 2740 11840 2746 11852
rect 3069 11849 3081 11852
rect 3115 11849 3127 11883
rect 3069 11843 3127 11849
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3878 11880 3884 11892
rect 3283 11852 3884 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 1949 11815 2007 11821
rect 1949 11812 1961 11815
rect 1912 11784 1961 11812
rect 1912 11772 1918 11784
rect 1949 11781 1961 11784
rect 1995 11781 2007 11815
rect 1949 11775 2007 11781
rect 2869 11815 2927 11821
rect 2869 11781 2881 11815
rect 2915 11812 2927 11815
rect 2958 11812 2964 11824
rect 2915 11784 2964 11812
rect 2915 11781 2927 11784
rect 2869 11775 2927 11781
rect 2958 11772 2964 11784
rect 3016 11772 3022 11824
rect 1578 11704 1584 11756
rect 1636 11704 1642 11756
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2096 11716 2237 11744
rect 2096 11704 2102 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3234 11744 3240 11756
rect 2547 11716 3240 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 3344 11753 3372 11852
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4982 11880 4988 11892
rect 4080 11852 4988 11880
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3602 11704 3608 11756
rect 3660 11704 3666 11756
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 4080 11753 4108 11852
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 5224 11852 5273 11880
rect 5224 11840 5230 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 6546 11840 6552 11892
rect 6604 11840 6610 11892
rect 7466 11880 7472 11892
rect 6840 11852 7472 11880
rect 4430 11772 4436 11824
rect 4488 11812 4494 11824
rect 4706 11812 4712 11824
rect 4488 11784 4712 11812
rect 4488 11772 4494 11784
rect 4706 11772 4712 11784
rect 4764 11812 4770 11824
rect 5077 11815 5135 11821
rect 5077 11812 5089 11815
rect 4764 11784 5089 11812
rect 4764 11772 4770 11784
rect 5077 11781 5089 11784
rect 5123 11781 5135 11815
rect 5994 11812 6000 11824
rect 5077 11775 5135 11781
rect 5460 11784 6000 11812
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3970 11676 3976 11688
rect 2639 11648 3976 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 4080 11608 4108 11707
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4338 11744 4344 11756
rect 4295 11716 4344 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4338 11704 4344 11716
rect 4396 11744 4402 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4396 11716 4813 11744
rect 4396 11704 4402 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 5460 11753 5488 11784
rect 5994 11772 6000 11784
rect 6052 11812 6058 11824
rect 6052 11784 6776 11812
rect 6052 11772 6058 11784
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5040 11716 5457 11744
rect 5040 11704 5046 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5534 11704 5540 11756
rect 5592 11704 5598 11756
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 6748 11753 6776 11784
rect 6840 11753 6868 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 7800 11852 8953 11880
rect 7800 11840 7806 11852
rect 8941 11849 8953 11852
rect 8987 11849 8999 11883
rect 8941 11843 8999 11849
rect 7285 11815 7343 11821
rect 7285 11781 7297 11815
rect 7331 11812 7343 11815
rect 7331 11784 8248 11812
rect 7331 11781 7343 11784
rect 7285 11775 7343 11781
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 6972 11716 7113 11744
rect 6972 11704 6978 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7190 11704 7196 11756
rect 7248 11704 7254 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 4172 11676 4200 11704
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 4172 11648 4721 11676
rect 4709 11645 4721 11648
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 7392 11676 7420 11707
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 7558 11704 7564 11756
rect 7616 11704 7622 11756
rect 7742 11704 7748 11756
rect 7800 11704 7806 11756
rect 8220 11753 8248 11784
rect 8294 11772 8300 11824
rect 8352 11812 8358 11824
rect 9217 11815 9275 11821
rect 8352 11784 8892 11812
rect 8352 11772 8358 11784
rect 8864 11753 8892 11784
rect 9217 11781 9229 11815
rect 9263 11812 9275 11815
rect 10226 11812 10232 11824
rect 9263 11784 10232 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 5767 11648 6040 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 4154 11608 4160 11620
rect 2924 11580 4016 11608
rect 4080 11580 4160 11608
rect 2924 11568 2930 11580
rect 1946 11500 1952 11552
rect 2004 11500 2010 11552
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3142 11540 3148 11552
rect 3099 11512 3148 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 3786 11500 3792 11552
rect 3844 11500 3850 11552
rect 3988 11540 4016 11580
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 4246 11568 4252 11620
rect 4304 11608 4310 11620
rect 4617 11611 4675 11617
rect 4617 11608 4629 11611
rect 4304 11580 4629 11608
rect 4304 11568 4310 11580
rect 4617 11577 4629 11580
rect 4663 11608 4675 11611
rect 5258 11608 5264 11620
rect 4663 11580 5264 11608
rect 4663 11577 4675 11580
rect 4617 11571 4675 11577
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 6012 11608 6040 11648
rect 6748 11648 7420 11676
rect 8297 11679 8355 11685
rect 6178 11608 6184 11620
rect 6012 11580 6184 11608
rect 4430 11540 4436 11552
rect 3988 11512 4436 11540
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4522 11500 4528 11552
rect 4580 11500 4586 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5166 11540 5172 11552
rect 4856 11512 5172 11540
rect 4856 11500 4862 11512
rect 5166 11500 5172 11512
rect 5224 11540 5230 11552
rect 6012 11540 6040 11580
rect 6178 11568 6184 11580
rect 6236 11608 6242 11620
rect 6748 11608 6776 11648
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8386 11676 8392 11688
rect 8343 11648 8392 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 9048 11676 9076 11707
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 8588 11648 9444 11676
rect 8588 11617 8616 11648
rect 6236 11580 6776 11608
rect 8573 11611 8631 11617
rect 6236 11568 6242 11580
rect 8573 11577 8585 11611
rect 8619 11577 8631 11611
rect 8573 11571 8631 11577
rect 8665 11611 8723 11617
rect 8665 11577 8677 11611
rect 8711 11577 8723 11611
rect 8665 11571 8723 11577
rect 5224 11512 6040 11540
rect 5224 11500 5230 11512
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7006 11540 7012 11552
rect 6696 11512 7012 11540
rect 6696 11500 6702 11512
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7926 11500 7932 11552
rect 7984 11500 7990 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 8680 11540 8708 11571
rect 9416 11549 9444 11648
rect 8168 11512 8708 11540
rect 9401 11543 9459 11549
rect 8168 11500 8174 11512
rect 9401 11509 9413 11543
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 9769 11543 9827 11549
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 9858 11540 9864 11552
rect 9815 11512 9864 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 1104 11450 10856 11472
rect 1104 11398 2169 11450
rect 2221 11398 2233 11450
rect 2285 11398 2297 11450
rect 2349 11398 2361 11450
rect 2413 11398 2425 11450
rect 2477 11398 4607 11450
rect 4659 11398 4671 11450
rect 4723 11398 4735 11450
rect 4787 11398 4799 11450
rect 4851 11398 4863 11450
rect 4915 11398 7045 11450
rect 7097 11398 7109 11450
rect 7161 11398 7173 11450
rect 7225 11398 7237 11450
rect 7289 11398 7301 11450
rect 7353 11398 9483 11450
rect 9535 11398 9547 11450
rect 9599 11398 9611 11450
rect 9663 11398 9675 11450
rect 9727 11398 9739 11450
rect 9791 11398 10856 11450
rect 1104 11376 10856 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2590 11336 2596 11348
rect 2455 11308 2596 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 3418 11336 3424 11348
rect 3375 11308 3424 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 4154 11336 4160 11348
rect 3559 11308 4160 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5040 11308 5181 11336
rect 5040 11296 5046 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 6362 11336 6368 11348
rect 5583 11308 6368 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7466 11336 7472 11348
rect 7331 11308 7472 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7466 11296 7472 11308
rect 7524 11336 7530 11348
rect 8018 11336 8024 11348
rect 7524 11308 8024 11336
rect 7524 11296 7530 11308
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9048 11308 9689 11336
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11237 1639 11271
rect 1581 11231 1639 11237
rect 2133 11271 2191 11277
rect 2133 11237 2145 11271
rect 2179 11268 2191 11271
rect 2314 11268 2320 11280
rect 2179 11240 2320 11268
rect 2179 11237 2191 11240
rect 2133 11231 2191 11237
rect 1596 11200 1624 11231
rect 2314 11228 2320 11240
rect 2372 11268 2378 11280
rect 3234 11268 3240 11280
rect 2372 11240 3240 11268
rect 2372 11228 2378 11240
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 3786 11228 3792 11280
rect 3844 11268 3850 11280
rect 4338 11268 4344 11280
rect 3844 11240 4344 11268
rect 3844 11228 3850 11240
rect 3988 11209 4016 11240
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 4798 11268 4804 11280
rect 4488 11240 4804 11268
rect 4488 11228 4494 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 5077 11271 5135 11277
rect 5077 11237 5089 11271
rect 5123 11268 5135 11271
rect 5123 11240 7052 11268
rect 5123 11237 5135 11240
rect 5077 11231 5135 11237
rect 3973 11203 4031 11209
rect 1596 11172 2360 11200
rect 842 11092 848 11144
rect 900 11132 906 11144
rect 1397 11135 1455 11141
rect 1397 11132 1409 11135
rect 900 11104 1409 11132
rect 900 11092 906 11104
rect 1397 11101 1409 11104
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1765 11135 1823 11141
rect 1765 11132 1777 11135
rect 1636 11104 1777 11132
rect 1636 11092 1642 11104
rect 1765 11101 1777 11104
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1912 11104 1961 11132
rect 1912 11092 1918 11104
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 2332 11132 2360 11172
rect 2516 11172 3280 11200
rect 2516 11132 2544 11172
rect 3252 11144 3280 11172
rect 3973 11169 3985 11203
rect 4019 11169 4031 11203
rect 4246 11200 4252 11212
rect 3973 11163 4031 11169
rect 4080 11172 4252 11200
rect 2332 11104 2544 11132
rect 1949 11095 2007 11101
rect 2590 11092 2596 11144
rect 2648 11132 2654 11144
rect 3053 11135 3111 11141
rect 3053 11132 3065 11135
rect 2648 11104 3065 11132
rect 2648 11092 2654 11104
rect 3053 11101 3065 11104
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 4080 11141 4108 11172
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4580 11172 5212 11200
rect 4580 11160 4586 11172
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4212 11104 4445 11132
rect 4212 11092 4218 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4614 11092 4620 11144
rect 4672 11092 4678 11144
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 2038 11024 2044 11076
rect 2096 11064 2102 11076
rect 2225 11067 2283 11073
rect 2225 11064 2237 11067
rect 2096 11036 2237 11064
rect 2096 11024 2102 11036
rect 2225 11033 2237 11036
rect 2271 11033 2283 11067
rect 2225 11027 2283 11033
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 2425 11067 2483 11073
rect 2425 11064 2437 11067
rect 2372 11036 2437 11064
rect 2372 11024 2378 11036
rect 2425 11033 2437 11036
rect 2471 11033 2483 11067
rect 2866 11064 2872 11076
rect 2425 11027 2483 11033
rect 2608 11036 2872 11064
rect 2608 11005 2636 11036
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 3160 11064 3188 11092
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 3160 11036 3341 11064
rect 3329 11033 3341 11036
rect 3375 11064 3387 11067
rect 3510 11064 3516 11076
rect 3375 11036 3516 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 4341 11067 4399 11073
rect 4341 11033 4353 11067
rect 4387 11064 4399 11067
rect 4522 11064 4528 11076
rect 4387 11036 4528 11064
rect 4387 11033 4399 11036
rect 4341 11027 4399 11033
rect 4522 11024 4528 11036
rect 4580 11064 4586 11076
rect 4724 11064 4752 11095
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 5184 11141 5212 11172
rect 5258 11160 5264 11212
rect 5316 11160 5322 11212
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6914 11200 6920 11212
rect 6319 11172 6920 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6546 11132 6552 11144
rect 6503 11104 6552 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 7024 11132 7052 11240
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8202 11268 8208 11280
rect 7984 11240 8208 11268
rect 7984 11228 7990 11240
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9048 11268 9076 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 9861 11339 9919 11345
rect 9861 11336 9873 11339
rect 9824 11308 9873 11336
rect 9824 11296 9830 11308
rect 9861 11305 9873 11308
rect 9907 11305 9919 11339
rect 9861 11299 9919 11305
rect 8956 11240 9076 11268
rect 9585 11271 9643 11277
rect 8956 11209 8984 11240
rect 9585 11237 9597 11271
rect 9631 11268 9643 11271
rect 10042 11268 10048 11280
rect 9631 11240 10048 11268
rect 9631 11237 9643 11240
rect 9585 11231 9643 11237
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10226 11228 10232 11280
rect 10284 11268 10290 11280
rect 10502 11268 10508 11280
rect 10284 11240 10508 11268
rect 10284 11228 10290 11240
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 8946 11203 9004 11209
rect 8946 11169 8958 11203
rect 8992 11169 9004 11203
rect 8946 11163 9004 11169
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9766 11200 9772 11212
rect 9180 11172 9772 11200
rect 9180 11160 9186 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 7024 11104 9045 11132
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9404 11135 9462 11141
rect 9404 11132 9416 11135
rect 9033 11095 9091 11101
rect 9140 11104 9416 11132
rect 4580 11036 4752 11064
rect 6641 11067 6699 11073
rect 4580 11024 4586 11036
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 6687 11036 7052 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 2593 10999 2651 11005
rect 2593 10965 2605 10999
rect 2639 10965 2651 10999
rect 2593 10959 2651 10965
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3145 10999 3203 11005
rect 3145 10996 3157 10999
rect 3016 10968 3157 10996
rect 3016 10956 3022 10968
rect 3145 10965 3157 10968
rect 3191 10996 3203 10999
rect 4062 10996 4068 11008
rect 3191 10968 4068 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 7024 10996 7052 11036
rect 7098 11024 7104 11076
rect 7156 11024 7162 11076
rect 7301 11067 7359 11073
rect 7301 11064 7313 11067
rect 7208 11036 7313 11064
rect 7208 10996 7236 11036
rect 7301 11033 7313 11036
rect 7347 11064 7359 11067
rect 7742 11064 7748 11076
rect 7347 11036 7748 11064
rect 7347 11033 7359 11036
rect 7301 11027 7359 11033
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 7024 10968 7236 10996
rect 7469 10999 7527 11005
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7558 10996 7564 11008
rect 7515 10968 7564 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7558 10956 7564 10968
rect 7616 10996 7622 11008
rect 7944 10996 7972 11027
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 9140 11064 9168 11104
rect 9404 11101 9416 11104
rect 9450 11101 9462 11135
rect 9404 11095 9462 11101
rect 8076 11036 9168 11064
rect 8076 11024 8082 11036
rect 9858 11024 9864 11076
rect 9916 11024 9922 11076
rect 7616 10968 7972 10996
rect 7616 10956 7622 10968
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 9088 10968 9413 10996
rect 9088 10956 9094 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 9401 10959 9459 10965
rect 1104 10906 10856 10928
rect 1104 10854 2829 10906
rect 2881 10854 2893 10906
rect 2945 10854 2957 10906
rect 3009 10854 3021 10906
rect 3073 10854 3085 10906
rect 3137 10854 5267 10906
rect 5319 10854 5331 10906
rect 5383 10854 5395 10906
rect 5447 10854 5459 10906
rect 5511 10854 5523 10906
rect 5575 10854 7705 10906
rect 7757 10854 7769 10906
rect 7821 10854 7833 10906
rect 7885 10854 7897 10906
rect 7949 10854 7961 10906
rect 8013 10854 10143 10906
rect 10195 10854 10207 10906
rect 10259 10854 10271 10906
rect 10323 10854 10335 10906
rect 10387 10854 10399 10906
rect 10451 10854 10856 10906
rect 1104 10832 10856 10854
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4672 10764 4813 10792
rect 4672 10752 4678 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 5258 10792 5264 10804
rect 4801 10755 4859 10761
rect 4908 10764 5264 10792
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1670 10616 1676 10668
rect 1728 10616 1734 10668
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 4908 10656 4936 10764
rect 5258 10752 5264 10764
rect 5316 10792 5322 10804
rect 5718 10792 5724 10804
rect 5316 10764 5724 10792
rect 5316 10752 5322 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5994 10792 6000 10804
rect 5828 10764 6000 10792
rect 5828 10724 5856 10764
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 9030 10792 9036 10804
rect 6328 10764 9036 10792
rect 6328 10752 6334 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10410 10752 10416 10804
rect 10468 10752 10474 10804
rect 7374 10724 7380 10736
rect 5736 10696 5856 10724
rect 6012 10696 7380 10724
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4908 10628 4997 10656
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5353 10659 5411 10665
rect 5215 10628 5304 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4212 10560 4353 10588
rect 4212 10548 4218 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 1946 10520 1952 10532
rect 1627 10492 1952 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 4617 10523 4675 10529
rect 4617 10489 4629 10523
rect 4663 10520 4675 10523
rect 4890 10520 4896 10532
rect 4663 10492 4896 10520
rect 4663 10489 4675 10492
rect 4617 10483 4675 10489
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 1854 10412 1860 10464
rect 1912 10412 1918 10464
rect 4338 10412 4344 10464
rect 4396 10412 4402 10464
rect 5092 10452 5120 10619
rect 5276 10520 5304 10628
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5368 10588 5396 10619
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 5736 10665 5764 10696
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 6012 10600 6040 10696
rect 7374 10684 7380 10696
rect 7432 10724 7438 10736
rect 7432 10696 8156 10724
rect 7432 10684 7438 10696
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6914 10656 6920 10668
rect 6135 10628 6920 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5368 10560 5549 10588
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 5994 10548 6000 10600
rect 6052 10548 6058 10600
rect 5442 10520 5448 10532
rect 5276 10492 5448 10520
rect 5442 10480 5448 10492
rect 5500 10520 5506 10532
rect 6104 10520 6132 10619
rect 6914 10616 6920 10628
rect 6972 10656 6978 10668
rect 7466 10656 7472 10668
rect 6972 10628 7472 10656
rect 6972 10616 6978 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8128 10665 8156 10696
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7616 10628 7849 10656
rect 7616 10616 7622 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 8018 10588 8024 10600
rect 6236 10560 8024 10588
rect 6236 10548 6242 10560
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8128 10588 8156 10619
rect 8202 10616 8208 10668
rect 8260 10616 8266 10668
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 10100 10628 10241 10656
rect 10100 10616 10106 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 8128 10560 8248 10588
rect 8220 10532 8248 10560
rect 5500 10492 6132 10520
rect 5500 10480 5506 10492
rect 8202 10480 8208 10532
rect 8260 10480 8266 10532
rect 5994 10452 6000 10464
rect 5092 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 7837 10455 7895 10461
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8938 10452 8944 10464
rect 7883 10424 8944 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 1104 10362 10856 10384
rect 1104 10310 2169 10362
rect 2221 10310 2233 10362
rect 2285 10310 2297 10362
rect 2349 10310 2361 10362
rect 2413 10310 2425 10362
rect 2477 10310 4607 10362
rect 4659 10310 4671 10362
rect 4723 10310 4735 10362
rect 4787 10310 4799 10362
rect 4851 10310 4863 10362
rect 4915 10310 7045 10362
rect 7097 10310 7109 10362
rect 7161 10310 7173 10362
rect 7225 10310 7237 10362
rect 7289 10310 7301 10362
rect 7353 10310 9483 10362
rect 9535 10310 9547 10362
rect 9599 10310 9611 10362
rect 9663 10310 9675 10362
rect 9727 10310 9739 10362
rect 9791 10310 10856 10362
rect 1104 10288 10856 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 3970 10248 3976 10260
rect 3016 10220 3976 10248
rect 3016 10208 3022 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5166 10248 5172 10260
rect 4939 10220 5172 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5810 10248 5816 10260
rect 5675 10220 5816 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 1854 10140 1860 10192
rect 1912 10180 1918 10192
rect 6546 10180 6552 10192
rect 1912 10152 6552 10180
rect 1912 10140 1918 10152
rect 2240 10053 2268 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 8754 10140 8760 10192
rect 8812 10180 8818 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 8812 10152 9229 10180
rect 8812 10140 8818 10152
rect 9217 10149 9229 10152
rect 9263 10149 9275 10183
rect 9217 10143 9275 10149
rect 3878 10112 3884 10124
rect 2792 10084 3884 10112
rect 2792 10053 2820 10084
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 5994 10112 6000 10124
rect 4028 10084 6000 10112
rect 4028 10072 4034 10084
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2866 10004 2872 10056
rect 2924 10004 2930 10056
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 1486 9936 1492 9988
rect 1544 9936 1550 9988
rect 1670 9936 1676 9988
rect 1728 9936 1734 9988
rect 2038 9936 2044 9988
rect 2096 9976 2102 9988
rect 2593 9979 2651 9985
rect 2593 9976 2605 9979
rect 2096 9948 2605 9976
rect 2096 9936 2102 9948
rect 2593 9945 2605 9948
rect 2639 9945 2651 9979
rect 2593 9939 2651 9945
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3068 9976 3096 10007
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 5368 10053 5396 10084
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 8938 10072 8944 10124
rect 8996 10072 9002 10124
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 3384 10016 4721 10044
rect 3384 10004 3390 10016
rect 4709 10013 4721 10016
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 5442 10004 5448 10056
rect 5500 10004 5506 10056
rect 2740 9948 3096 9976
rect 5629 9979 5687 9985
rect 2740 9936 2746 9948
rect 5629 9945 5641 9979
rect 5675 9976 5687 9979
rect 5994 9976 6000 9988
rect 5675 9948 6000 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 1912 9880 2421 9908
rect 1912 9868 1918 9880
rect 2409 9877 2421 9880
rect 2455 9908 2467 9911
rect 2866 9908 2872 9920
rect 2455 9880 2872 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2866 9868 2872 9880
rect 2924 9908 2930 9920
rect 3510 9908 3516 9920
rect 2924 9880 3516 9908
rect 2924 9868 2930 9880
rect 3510 9868 3516 9880
rect 3568 9908 3574 9920
rect 6638 9908 6644 9920
rect 3568 9880 6644 9908
rect 3568 9868 3574 9880
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 9401 9911 9459 9917
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9674 9908 9680 9920
rect 9447 9880 9680 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 1104 9818 10856 9840
rect 1104 9766 2829 9818
rect 2881 9766 2893 9818
rect 2945 9766 2957 9818
rect 3009 9766 3021 9818
rect 3073 9766 3085 9818
rect 3137 9766 5267 9818
rect 5319 9766 5331 9818
rect 5383 9766 5395 9818
rect 5447 9766 5459 9818
rect 5511 9766 5523 9818
rect 5575 9766 7705 9818
rect 7757 9766 7769 9818
rect 7821 9766 7833 9818
rect 7885 9766 7897 9818
rect 7949 9766 7961 9818
rect 8013 9766 10143 9818
rect 10195 9766 10207 9818
rect 10259 9766 10271 9818
rect 10323 9766 10335 9818
rect 10387 9766 10399 9818
rect 10451 9766 10856 9818
rect 1104 9744 10856 9766
rect 1762 9664 1768 9716
rect 1820 9704 1826 9716
rect 2590 9704 2596 9716
rect 1820 9676 2596 9704
rect 1820 9664 1826 9676
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3970 9704 3976 9716
rect 3283 9676 3976 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 2774 9636 2780 9648
rect 1412 9608 2780 9636
rect 1412 9577 1440 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 3252 9636 3280 9667
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 4154 9664 4160 9716
rect 4212 9664 4218 9716
rect 4062 9636 4068 9648
rect 2884 9608 3280 9636
rect 3344 9608 4068 9636
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 1854 9568 1860 9580
rect 1535 9540 1860 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2884 9568 2912 9608
rect 2593 9531 2651 9537
rect 2746 9540 2912 9568
rect 3053 9571 3111 9577
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 1762 9500 1768 9512
rect 1719 9472 1768 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9469 2559 9503
rect 2608 9500 2636 9531
rect 2746 9500 2774 9540
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3234 9568 3240 9580
rect 3099 9540 3240 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 2608 9472 2774 9500
rect 2501 9463 2559 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 2516 9432 2544 9463
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3344 9500 3372 9608
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 6546 9596 6552 9648
rect 6604 9596 6610 9648
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 3786 9528 3792 9580
rect 3844 9528 3850 9580
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6236 9540 6653 9568
rect 6236 9528 6242 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 3200 9472 3372 9500
rect 3200 9460 3206 9472
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4982 9500 4988 9512
rect 4028 9472 4988 9500
rect 4028 9460 4034 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6748 9500 6776 9599
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8168 9608 9628 9636
rect 8168 9596 8174 9608
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 8754 9528 8760 9580
rect 8812 9528 8818 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9048 9540 9505 9568
rect 6144 9472 6776 9500
rect 6144 9460 6150 9472
rect 1627 9404 2544 9432
rect 2961 9435 3019 9441
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 2961 9401 2973 9435
rect 3007 9432 3019 9435
rect 3896 9432 3924 9460
rect 3007 9404 3924 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 5350 9432 5356 9444
rect 4120 9404 5356 9432
rect 4120 9392 4126 9404
rect 5350 9392 5356 9404
rect 5408 9432 5414 9444
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 5408 9404 6377 9432
rect 5408 9392 5414 9404
rect 6365 9401 6377 9404
rect 6411 9432 6423 9435
rect 6840 9432 6868 9528
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 8018 9500 8024 9512
rect 6972 9472 8024 9500
rect 6972 9460 6978 9472
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 8938 9500 8944 9512
rect 8895 9472 8944 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 6411 9404 6868 9432
rect 6411 9401 6423 9404
rect 6365 9395 6423 9401
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 9048 9432 9076 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9398 9500 9404 9512
rect 9140 9472 9404 9500
rect 9140 9441 9168 9472
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 8352 9404 9076 9432
rect 9125 9435 9183 9441
rect 8352 9392 8358 9404
rect 9125 9401 9137 9435
rect 9171 9401 9183 9435
rect 9508 9432 9536 9531
rect 9600 9509 9628 9608
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 9861 9531 9919 9537
rect 9968 9540 10057 9568
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9876 9500 9904 9531
rect 9631 9472 9904 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 9968 9432 9996 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 9508 9404 9996 9432
rect 9125 9395 9183 9401
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 3142 9364 3148 9376
rect 2271 9336 3148 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 6270 9364 6276 9376
rect 3292 9336 6276 9364
rect 3292 9324 3298 9336
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6914 9324 6920 9376
rect 6972 9324 6978 9376
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9364 9336 9965 9364
rect 9364 9324 9370 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2004 9132 2697 9160
rect 2004 9120 2010 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3234 9160 3240 9172
rect 2823 9132 3240 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2700 9024 2728 9123
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3936 9132 4077 9160
rect 3936 9120 3942 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 6457 9163 6515 9169
rect 4755 9132 6224 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 3510 9092 3516 9104
rect 2915 9064 3516 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 2700 8996 3188 9024
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1544 8928 1685 8956
rect 1544 8916 1550 8928
rect 1673 8925 1685 8928
rect 1719 8956 1731 8959
rect 2498 8956 2504 8968
rect 1719 8928 2504 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 3160 8965 3188 8996
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 4724 9024 4752 9123
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 6086 9092 6092 9104
rect 5592 9064 6092 9092
rect 5592 9052 5598 9064
rect 6086 9052 6092 9064
rect 6144 9052 6150 9104
rect 6196 9092 6224 9132
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 7006 9160 7012 9172
rect 6503 9132 7012 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8754 9160 8760 9172
rect 7975 9132 8760 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 6730 9092 6736 9104
rect 6196 9064 6736 9092
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 6914 9052 6920 9104
rect 6972 9052 6978 9104
rect 10413 9095 10471 9101
rect 10413 9092 10425 9095
rect 9968 9064 10425 9092
rect 3844 8996 4752 9024
rect 5629 9027 5687 9033
rect 3844 8984 3850 8996
rect 3988 8965 4016 8996
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 6748 9024 6776 9052
rect 5675 8996 6408 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8956 4583 8959
rect 5718 8956 5724 8968
rect 5776 8965 5782 8968
rect 4571 8928 5724 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 4540 8888 4568 8919
rect 5718 8916 5724 8928
rect 5776 8919 5784 8965
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8950 5963 8959
rect 5951 8925 6045 8950
rect 5905 8922 6045 8925
rect 5905 8919 5963 8922
rect 5776 8916 5782 8919
rect 1912 8860 4568 8888
rect 1912 8848 1918 8860
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8857 5687 8891
rect 5629 8851 5687 8857
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 2096 8792 2329 8820
rect 2096 8780 2102 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2317 8783 2375 8789
rect 3329 8823 3387 8829
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 4062 8820 4068 8832
rect 3375 8792 4068 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 4396 8792 4445 8820
rect 4396 8780 4402 8792
rect 4433 8789 4445 8792
rect 4479 8789 4491 8823
rect 5644 8820 5672 8851
rect 6017 8820 6045 8922
rect 6178 8916 6184 8968
rect 6236 8916 6242 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6086 8848 6092 8900
rect 6144 8848 6150 8900
rect 6380 8888 6408 8996
rect 6564 8996 6776 9024
rect 6564 8965 6592 8996
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 6696 8928 6745 8956
rect 6696 8916 6702 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7432 8928 7665 8956
rect 7432 8916 7438 8928
rect 7653 8925 7665 8928
rect 7699 8956 7711 8959
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7699 8928 7757 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 6917 8891 6975 8897
rect 6917 8888 6929 8891
rect 6380 8860 6929 8888
rect 6917 8857 6929 8860
rect 6963 8888 6975 8891
rect 7098 8888 7104 8900
rect 6963 8860 7104 8888
rect 6963 8857 6975 8860
rect 6917 8851 6975 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7340 8860 7512 8888
rect 7340 8848 7346 8860
rect 6546 8820 6552 8832
rect 5644 8792 6552 8820
rect 4433 8783 4491 8789
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7484 8829 7512 8860
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 7944 8888 7972 8919
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9968 8965 9996 9064
rect 10413 9061 10425 9064
rect 10459 9061 10471 9095
rect 10413 9055 10471 9061
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10100 8996 10241 9024
rect 10100 8984 10106 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9692 8928 9965 8956
rect 7616 8860 7972 8888
rect 8036 8860 8248 8888
rect 7616 8848 7622 8860
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 7248 8792 7389 8820
rect 7248 8780 7254 8792
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 7469 8823 7527 8829
rect 7469 8789 7481 8823
rect 7515 8820 7527 8823
rect 8036 8820 8064 8860
rect 8220 8832 8248 8860
rect 7515 8792 8064 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 8110 8780 8116 8832
rect 8168 8780 8174 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 9692 8829 9720 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10502 8956 10508 8968
rect 10183 8928 10508 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 9769 8891 9827 8897
rect 9769 8857 9781 8891
rect 9815 8888 9827 8891
rect 10042 8888 10048 8900
rect 9815 8860 10048 8888
rect 9815 8857 9827 8860
rect 9769 8851 9827 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8789 9735 8823
rect 9677 8783 9735 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 9916 8792 10241 8820
rect 9916 8780 9922 8792
rect 10229 8789 10241 8792
rect 10275 8789 10287 8823
rect 10229 8783 10287 8789
rect 1104 8730 10856 8752
rect 1104 8678 2829 8730
rect 2881 8678 2893 8730
rect 2945 8678 2957 8730
rect 3009 8678 3021 8730
rect 3073 8678 3085 8730
rect 3137 8678 5267 8730
rect 5319 8678 5331 8730
rect 5383 8678 5395 8730
rect 5447 8678 5459 8730
rect 5511 8678 5523 8730
rect 5575 8678 7705 8730
rect 7757 8678 7769 8730
rect 7821 8678 7833 8730
rect 7885 8678 7897 8730
rect 7949 8678 7961 8730
rect 8013 8678 10143 8730
rect 10195 8678 10207 8730
rect 10259 8678 10271 8730
rect 10323 8678 10335 8730
rect 10387 8678 10399 8730
rect 10451 8678 10856 8730
rect 1104 8656 10856 8678
rect 7282 8576 7288 8628
rect 7340 8576 7346 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7558 8616 7564 8628
rect 7515 8588 7564 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 10413 8619 10471 8625
rect 8260 8588 8616 8616
rect 8260 8576 8266 8588
rect 6089 8551 6147 8557
rect 4264 8520 5120 8548
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 4264 8489 4292 8520
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3292 8452 4261 8480
rect 3292 8440 3298 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8478 4583 8483
rect 4614 8478 4620 8492
rect 4571 8450 4620 8478
rect 4571 8449 4583 8450
rect 4525 8443 4583 8449
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 1762 8412 1768 8424
rect 1719 8384 1768 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 4448 8412 4476 8443
rect 4614 8440 4620 8450
rect 4672 8440 4678 8492
rect 5092 8489 5120 8520
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6454 8548 6460 8560
rect 6135 8520 6460 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 8588 8557 8616 8588
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10870 8616 10876 8628
rect 10459 8588 10876 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 8357 8551 8415 8557
rect 8357 8548 8369 8551
rect 6696 8520 8369 8548
rect 6696 8508 6702 8520
rect 8357 8517 8369 8520
rect 8403 8517 8415 8551
rect 8357 8511 8415 8517
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8517 8631 8551
rect 8573 8511 8631 8517
rect 8680 8520 9536 8548
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5994 8480 6000 8492
rect 5307 8452 6000 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5276 8412 5304 8443
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6270 8480 6276 8492
rect 6227 8452 6276 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6779 8452 7236 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 4448 8384 5304 8412
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8412 6975 8415
rect 7098 8412 7104 8424
rect 6963 8384 7104 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7208 8412 7236 8452
rect 7282 8440 7288 8492
rect 7340 8489 7346 8492
rect 7340 8483 7402 8489
rect 7340 8449 7356 8483
rect 7390 8480 7402 8483
rect 7466 8480 7472 8492
rect 7390 8452 7472 8480
rect 7390 8449 7402 8452
rect 7340 8443 7402 8449
rect 7340 8440 7346 8443
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7791 8452 8248 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 7208 8384 7849 8412
rect 7837 8381 7849 8384
rect 7883 8412 7895 8415
rect 8018 8412 8024 8424
rect 7883 8384 8024 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 4614 8344 4620 8356
rect 4356 8316 4620 8344
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4356 8285 4384 8316
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 5077 8347 5135 8353
rect 5077 8344 5089 8347
rect 4816 8316 5089 8344
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 4212 8248 4353 8276
rect 4212 8236 4218 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 4341 8239 4399 8245
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4816 8285 4844 8316
rect 5077 8313 5089 8316
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 6730 8344 6736 8356
rect 6503 8316 6736 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 8110 8304 8116 8356
rect 8168 8304 8174 8356
rect 8220 8353 8248 8452
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8313 8263 8347
rect 8680 8344 8708 8520
rect 8938 8440 8944 8492
rect 8996 8440 9002 8492
rect 9508 8489 9536 8520
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 9263 8452 9321 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 9858 8480 9864 8492
rect 9815 8452 9864 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 8205 8307 8263 8313
rect 8312 8316 8708 8344
rect 4801 8279 4859 8285
rect 4801 8276 4813 8279
rect 4488 8248 4813 8276
rect 4488 8236 4494 8248
rect 4801 8245 4813 8248
rect 4847 8245 4859 8279
rect 4801 8239 4859 8245
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 8312 8276 8340 8316
rect 5684 8248 8340 8276
rect 5684 8236 5690 8248
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 9048 8276 9076 8443
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10042 8480 10048 8492
rect 9999 8452 10048 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10244 8412 10272 8443
rect 9232 8384 10272 8412
rect 9232 8353 9260 8384
rect 9217 8347 9275 8353
rect 9217 8313 9229 8347
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 8444 8248 9076 8276
rect 8444 8236 8450 8248
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1728 8044 2176 8072
rect 1728 8032 1734 8044
rect 2038 7964 2044 8016
rect 2096 7964 2102 8016
rect 2148 8013 2176 8044
rect 2590 8032 2596 8084
rect 2648 8072 2654 8084
rect 2648 8044 3004 8072
rect 2648 8032 2654 8044
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 8004 2191 8007
rect 2682 8004 2688 8016
rect 2179 7976 2688 8004
rect 2179 7973 2191 7976
rect 2133 7967 2191 7973
rect 2682 7964 2688 7976
rect 2740 8004 2746 8016
rect 2740 7976 2912 8004
rect 2740 7964 2746 7976
rect 2056 7936 2084 7964
rect 2056 7908 2728 7936
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2498 7868 2504 7880
rect 2271 7840 2504 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 1964 7800 1992 7831
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2700 7877 2728 7908
rect 2884 7877 2912 7976
rect 2976 7877 3004 8044
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 5074 8072 5080 8084
rect 4764 8044 5080 8072
rect 4764 8032 4770 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5626 8072 5632 8084
rect 5491 8044 5632 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6512 8044 6745 8072
rect 6512 8032 6518 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 7208 8044 7880 8072
rect 4614 8004 4620 8016
rect 4356 7976 4620 8004
rect 4356 7948 4384 7976
rect 4614 7964 4620 7976
rect 4672 8004 4678 8016
rect 4672 7976 4844 8004
rect 4672 7964 4678 7976
rect 4338 7896 4344 7948
rect 4396 7896 4402 7948
rect 4430 7896 4436 7948
rect 4488 7896 4494 7948
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 4816 7945 4844 7976
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 5994 7936 6000 7948
rect 5276 7908 6000 7936
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4522 7868 4528 7880
rect 4295 7840 4528 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 5276 7877 5304 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6638 7896 6644 7948
rect 6696 7896 6702 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7208 7945 7236 8044
rect 7852 8013 7880 8044
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6880 7908 7205 7936
rect 6880 7896 6886 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7374 7936 7380 7948
rect 7331 7908 7380 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7374 7896 7380 7908
rect 7432 7936 7438 7948
rect 7432 7908 7788 7936
rect 7432 7896 7438 7908
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 2590 7800 2596 7812
rect 1964 7772 2596 7800
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 4540 7800 4568 7828
rect 4908 7800 4936 7831
rect 5074 7800 5080 7812
rect 4540 7772 5080 7800
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 5460 7800 5488 7831
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 5184 7772 5488 7800
rect 7101 7803 7159 7809
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 2498 7692 2504 7744
rect 2556 7692 2562 7744
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 5184 7741 5212 7772
rect 7101 7769 7113 7803
rect 7147 7800 7159 7803
rect 7484 7800 7512 7831
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7760 7877 7788 7908
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7616 7840 7665 7868
rect 7616 7828 7622 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 8021 7803 8079 7809
rect 8021 7800 8033 7803
rect 7147 7772 8033 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8021 7769 8033 7772
rect 8067 7769 8079 7803
rect 8021 7763 8079 7769
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3936 7704 3985 7732
rect 3936 7692 3942 7704
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 7524 7704 7757 7732
rect 7524 7692 7530 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 7745 7695 7803 7701
rect 1104 7642 10856 7664
rect 1104 7590 2829 7642
rect 2881 7590 2893 7642
rect 2945 7590 2957 7642
rect 3009 7590 3021 7642
rect 3073 7590 3085 7642
rect 3137 7590 5267 7642
rect 5319 7590 5331 7642
rect 5383 7590 5395 7642
rect 5447 7590 5459 7642
rect 5511 7590 5523 7642
rect 5575 7590 7705 7642
rect 7757 7590 7769 7642
rect 7821 7590 7833 7642
rect 7885 7590 7897 7642
rect 7949 7590 7961 7642
rect 8013 7590 10143 7642
rect 10195 7590 10207 7642
rect 10259 7590 10271 7642
rect 10323 7590 10335 7642
rect 10387 7590 10399 7642
rect 10451 7590 10856 7642
rect 1104 7568 10856 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 2317 7531 2375 7537
rect 1452 7500 1808 7528
rect 1452 7488 1458 7500
rect 1780 7472 1808 7500
rect 2317 7497 2329 7531
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 1820 7432 2268 7460
rect 1820 7420 1826 7432
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1728 7364 1961 7392
rect 1728 7352 1734 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2038 7284 2044 7336
rect 2096 7284 2102 7336
rect 2240 7324 2268 7432
rect 2332 7392 2360 7491
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 4982 7488 4988 7540
rect 5040 7488 5046 7540
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 4448 7460 4476 7488
rect 5000 7460 5028 7488
rect 5261 7463 5319 7469
rect 5261 7460 5273 7463
rect 2648 7432 2728 7460
rect 4448 7432 4752 7460
rect 5000 7432 5273 7460
rect 2648 7420 2654 7432
rect 2700 7401 2728 7432
rect 2685 7395 2743 7401
rect 2332 7364 2636 7392
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 2240 7296 2421 7324
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2608 7324 2636 7364
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 3234 7324 3240 7336
rect 2608 7296 3240 7324
rect 2409 7287 2467 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 4080 7324 4108 7355
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 4614 7352 4620 7404
rect 4672 7352 4678 7404
rect 4724 7401 4752 7432
rect 5261 7429 5273 7432
rect 5307 7429 5319 7463
rect 5261 7423 5319 7429
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 4908 7324 4936 7352
rect 5092 7324 5120 7355
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 4080 7296 4936 7324
rect 5000 7296 5120 7324
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 3973 7259 4031 7265
rect 1627 7228 2636 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2406 7188 2412 7200
rect 2096 7160 2412 7188
rect 2096 7148 2102 7160
rect 2406 7148 2412 7160
rect 2464 7188 2470 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 2464 7160 2513 7188
rect 2464 7148 2470 7160
rect 2501 7157 2513 7160
rect 2547 7157 2559 7191
rect 2608 7188 2636 7228
rect 3973 7225 3985 7259
rect 4019 7256 4031 7259
rect 4430 7256 4436 7268
rect 4019 7228 4436 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 5000 7256 5028 7296
rect 4672 7228 5028 7256
rect 5261 7259 5319 7265
rect 4672 7216 4678 7228
rect 5261 7225 5273 7259
rect 5307 7256 5319 7259
rect 5994 7256 6000 7268
rect 5307 7228 6000 7256
rect 5307 7225 5319 7228
rect 5261 7219 5319 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 2774 7188 2780 7200
rect 2608 7160 2780 7188
rect 2501 7151 2559 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 4154 7188 4160 7200
rect 2915 7160 4160 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4246 7148 4252 7200
rect 4304 7148 4310 7200
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5074 7188 5080 7200
rect 4764 7160 5080 7188
rect 4764 7148 4770 7160
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 5629 6987 5687 6993
rect 2832 6956 5580 6984
rect 2832 6944 2838 6956
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6885 2007 6919
rect 1949 6879 2007 6885
rect 1964 6848 1992 6879
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2682 6916 2688 6928
rect 2464 6888 2688 6916
rect 2464 6876 2470 6888
rect 2682 6876 2688 6888
rect 2740 6916 2746 6928
rect 2740 6888 3372 6916
rect 2740 6876 2746 6888
rect 3237 6851 3295 6857
rect 1964 6820 3096 6848
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1578 6740 1584 6792
rect 1636 6740 1642 6792
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1762 6780 1768 6792
rect 1719 6752 1768 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1762 6740 1768 6752
rect 1820 6780 1826 6792
rect 1820 6752 2084 6780
rect 1820 6740 1826 6752
rect 1596 6712 1624 6740
rect 1946 6712 1952 6724
rect 1596 6684 1952 6712
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2056 6712 2084 6752
rect 2222 6740 2228 6792
rect 2280 6740 2286 6792
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 2317 6715 2375 6721
rect 2317 6712 2329 6715
rect 2056 6684 2329 6712
rect 2317 6681 2329 6684
rect 2363 6681 2375 6715
rect 2608 6712 2636 6743
rect 2682 6740 2688 6792
rect 2740 6740 2746 6792
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3068 6789 3096 6820
rect 3237 6817 3249 6851
rect 3283 6817 3295 6851
rect 3237 6811 3295 6817
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2608 6684 2789 6712
rect 2317 6675 2375 6681
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 3252 6712 3280 6811
rect 3344 6789 3372 6888
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4614 6916 4620 6928
rect 4212 6888 4620 6916
rect 4212 6876 4218 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 5552 6916 5580 6956
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5718 6984 5724 6996
rect 5675 6956 5724 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 9769 6987 9827 6993
rect 9769 6953 9781 6987
rect 9815 6984 9827 6987
rect 10226 6984 10232 6996
rect 9815 6956 10232 6984
rect 9815 6953 9827 6956
rect 9769 6947 9827 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 6638 6916 6644 6928
rect 5552 6888 6644 6916
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 7208 6888 8340 6916
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 4028 6820 4353 6848
rect 4028 6808 4034 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4430 6808 4436 6860
rect 4488 6808 4494 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 4632 6820 5028 6848
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 3418 6712 3424 6724
rect 3252 6684 3424 6712
rect 2777 6675 2835 6681
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 1578 6604 1584 6656
rect 1636 6604 1642 6656
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 1765 6647 1823 6653
rect 1765 6644 1777 6647
rect 1728 6616 1777 6644
rect 1728 6604 1734 6616
rect 1765 6613 1777 6616
rect 1811 6613 1823 6647
rect 1765 6607 1823 6613
rect 2041 6647 2099 6653
rect 2041 6613 2053 6647
rect 2087 6644 2099 6647
rect 4172 6644 4200 6743
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4632 6780 4660 6820
rect 4448 6752 4660 6780
rect 4448 6724 4476 6752
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 5000 6789 5028 6820
rect 5092 6820 5733 6848
rect 5092 6789 5120 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 5721 6811 5779 6817
rect 5828 6820 6193 6848
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5626 6780 5632 6792
rect 5552 6752 5632 6780
rect 4430 6672 4436 6724
rect 4488 6672 4494 6724
rect 4632 6684 5212 6712
rect 4632 6653 4660 6684
rect 2087 6616 4200 6644
rect 4617 6647 4675 6653
rect 2087 6613 2099 6616
rect 2041 6607 2099 6613
rect 4617 6613 4629 6647
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 4798 6604 4804 6656
rect 4856 6604 4862 6656
rect 5184 6644 5212 6684
rect 5258 6672 5264 6724
rect 5316 6672 5322 6724
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5552 6712 5580 6752
rect 5626 6740 5632 6752
rect 5684 6780 5690 6792
rect 5828 6780 5856 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 5684 6752 5856 6780
rect 5684 6740 5690 6752
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 7208 6780 7236 6888
rect 7300 6820 7604 6848
rect 7300 6789 7328 6820
rect 7576 6792 7604 6820
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 8168 6820 8217 6848
rect 8168 6808 8174 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8312 6848 8340 6888
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9490 6916 9496 6928
rect 9088 6888 9496 6916
rect 9088 6876 9094 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 9861 6919 9919 6925
rect 9861 6885 9873 6919
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 8312 6820 9628 6848
rect 8205 6811 8263 6817
rect 6420 6752 7236 6780
rect 7285 6783 7343 6789
rect 6420 6740 6426 6752
rect 7285 6749 7297 6783
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7616 6752 7941 6780
rect 7616 6740 7622 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8386 6780 8392 6792
rect 8067 6752 8392 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9214 6780 9220 6792
rect 9171 6752 9220 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9600 6789 9628 6820
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9876 6780 9904 6879
rect 9815 6752 9904 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10100 6752 10149 6780
rect 10100 6740 10106 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 5399 6684 5580 6712
rect 5920 6712 5948 6740
rect 6730 6712 6736 6724
rect 5920 6684 6736 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 9861 6715 9919 6721
rect 9861 6712 9873 6715
rect 7300 6684 9873 6712
rect 7300 6644 7328 6684
rect 9861 6681 9873 6684
rect 9907 6681 9919 6715
rect 9861 6675 9919 6681
rect 5184 6616 7328 6644
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7466 6644 7472 6656
rect 7423 6616 7472 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 8202 6604 8208 6656
rect 8260 6604 8266 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8720 6616 8953 6644
rect 8720 6604 8726 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 9824 6616 10057 6644
rect 9824 6604 9830 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 1104 6554 10856 6576
rect 1104 6502 2829 6554
rect 2881 6502 2893 6554
rect 2945 6502 2957 6554
rect 3009 6502 3021 6554
rect 3073 6502 3085 6554
rect 3137 6502 5267 6554
rect 5319 6502 5331 6554
rect 5383 6502 5395 6554
rect 5447 6502 5459 6554
rect 5511 6502 5523 6554
rect 5575 6502 7705 6554
rect 7757 6502 7769 6554
rect 7821 6502 7833 6554
rect 7885 6502 7897 6554
rect 7949 6502 7961 6554
rect 8013 6502 10143 6554
rect 10195 6502 10207 6554
rect 10259 6502 10271 6554
rect 10323 6502 10335 6554
rect 10387 6502 10399 6554
rect 10451 6502 10856 6554
rect 1104 6480 10856 6502
rect 1578 6400 1584 6452
rect 1636 6440 1642 6452
rect 3326 6440 3332 6452
rect 1636 6412 3332 6440
rect 1636 6400 1642 6412
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 4706 6440 4712 6452
rect 3651 6412 4712 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5868 6412 5917 6440
rect 5868 6400 5874 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 6362 6440 6368 6452
rect 5905 6403 5963 6409
rect 6012 6412 6368 6440
rect 1946 6372 1952 6384
rect 1596 6344 1952 6372
rect 1596 6316 1624 6344
rect 1946 6332 1952 6344
rect 2004 6332 2010 6384
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 3789 6375 3847 6381
rect 3292 6344 3740 6372
rect 3292 6332 3298 6344
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 3418 6304 3424 6316
rect 1820 6276 3424 6304
rect 1820 6264 1826 6276
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3712 6313 3740 6344
rect 3789 6341 3801 6375
rect 3835 6372 3847 6375
rect 4154 6372 4160 6384
rect 3835 6344 4160 6372
rect 3835 6341 3847 6344
rect 3789 6335 3847 6341
rect 4154 6332 4160 6344
rect 4212 6372 4218 6384
rect 4890 6372 4896 6384
rect 4212 6344 4896 6372
rect 4212 6332 4218 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 6012 6372 6040 6412
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8221 6443 8279 6449
rect 8221 6440 8233 6443
rect 7524 6412 8233 6440
rect 7524 6400 7530 6412
rect 8221 6409 8233 6412
rect 8267 6409 8279 6443
rect 8221 6403 8279 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8444 6412 8616 6440
rect 8444 6400 8450 6412
rect 5000 6344 6040 6372
rect 7193 6375 7251 6381
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 5000 6304 5028 6344
rect 7193 6341 7205 6375
rect 7239 6372 7251 6375
rect 7239 6344 7604 6372
rect 7239 6341 7251 6344
rect 7193 6335 7251 6341
rect 3927 6276 5028 6304
rect 5813 6307 5871 6313
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2222 6236 2228 6248
rect 2004 6208 2228 6236
rect 2004 6196 2010 6208
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 3436 6236 3464 6264
rect 3896 6236 3924 6267
rect 3436 6208 3924 6236
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 5626 6236 5632 6248
rect 4120 6208 5632 6236
rect 4120 6196 4126 6208
rect 5626 6196 5632 6208
rect 5684 6236 5690 6248
rect 5828 6236 5856 6267
rect 6086 6264 6092 6316
rect 6144 6264 6150 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6236 6276 6377 6304
rect 6236 6264 6242 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7116 6236 7144 6267
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7576 6313 7604 6344
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 8021 6375 8079 6381
rect 8021 6372 8033 6375
rect 7892 6344 8033 6372
rect 7892 6332 7898 6344
rect 8021 6341 8033 6344
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 8110 6264 8116 6316
rect 8168 6304 8174 6316
rect 8588 6313 8616 6412
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8168 6276 8493 6304
rect 8168 6264 8174 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8996 6276 9045 6304
rect 8996 6264 9002 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9033 6267 9091 6273
rect 9416 6276 9689 6304
rect 7374 6236 7380 6248
rect 5684 6208 7380 6236
rect 5684 6196 5690 6208
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7466 6196 7472 6248
rect 7524 6196 7530 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 7708 6208 8769 6236
rect 7708 6196 7714 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6089 6171 6147 6177
rect 6089 6168 6101 6171
rect 6052 6140 6101 6168
rect 6052 6128 6058 6140
rect 6089 6137 6101 6140
rect 6135 6137 6147 6171
rect 6089 6131 6147 6137
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 6549 6171 6607 6177
rect 6549 6168 6561 6171
rect 6328 6140 6561 6168
rect 6328 6128 6334 6140
rect 6549 6137 6561 6140
rect 6595 6137 6607 6171
rect 6549 6131 6607 6137
rect 6822 6128 6828 6180
rect 6880 6168 6886 6180
rect 7282 6168 7288 6180
rect 6880 6140 7288 6168
rect 6880 6128 6886 6140
rect 7282 6128 7288 6140
rect 7340 6168 7346 6180
rect 7834 6168 7840 6180
rect 7340 6140 7840 6168
rect 7340 6128 7346 6140
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 7929 6171 7987 6177
rect 7929 6137 7941 6171
rect 7975 6168 7987 6171
rect 9048 6168 9076 6267
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9214 6236 9220 6248
rect 9171 6208 9220 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9416 6245 9444 6276
rect 9677 6273 9689 6276
rect 9723 6304 9735 6307
rect 9858 6304 9864 6316
rect 9723 6276 9864 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 9950 6236 9956 6248
rect 9815 6208 9956 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 7975 6140 9076 6168
rect 7975 6137 7987 6140
rect 7929 6131 7987 6137
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 4338 6100 4344 6112
rect 2648 6072 4344 6100
rect 2648 6060 2654 6072
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7432 6072 8217 6100
rect 7432 6060 7438 6072
rect 8205 6069 8217 6072
rect 8251 6100 8263 6103
rect 8294 6100 8300 6112
rect 8251 6072 8300 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 6822 5896 6828 5908
rect 1627 5868 6828 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 7432 5868 7573 5896
rect 7432 5856 7438 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 5905 5831 5963 5837
rect 5905 5797 5917 5831
rect 5951 5828 5963 5831
rect 5994 5828 6000 5840
rect 5951 5800 6000 5828
rect 5951 5797 5963 5800
rect 5905 5791 5963 5797
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 7742 5788 7748 5840
rect 7800 5788 7806 5840
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 7926 5828 7932 5840
rect 7883 5800 7932 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8260 5800 9229 5828
rect 8260 5788 8266 5800
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5760 2191 5763
rect 2498 5760 2504 5772
rect 2179 5732 2504 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 7466 5760 7472 5772
rect 6144 5732 7472 5760
rect 6144 5720 6150 5732
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8496 5732 8953 5760
rect 8496 5704 8524 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1544 5664 2053 5692
rect 1544 5652 1550 5664
rect 2041 5661 2053 5664
rect 2087 5692 2099 5695
rect 2222 5692 2228 5704
rect 2087 5664 2228 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 4396 5664 5733 5692
rect 4396 5652 4402 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 6972 5664 7849 5692
rect 6972 5652 6978 5664
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 7576 5633 7604 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8294 5692 8300 5704
rect 8159 5664 8300 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8478 5652 8484 5704
rect 8536 5652 8542 5704
rect 8662 5652 8668 5704
rect 8720 5652 8726 5704
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 9048 5692 9076 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 8803 5664 9076 5692
rect 9493 5695 9551 5701
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 7377 5627 7435 5633
rect 7377 5624 7389 5627
rect 6328 5596 7389 5624
rect 6328 5584 6334 5596
rect 7377 5593 7389 5596
rect 7423 5593 7435 5627
rect 7576 5627 7635 5633
rect 7576 5596 7589 5627
rect 7377 5587 7435 5593
rect 7577 5593 7589 5596
rect 7623 5593 7635 5627
rect 8680 5624 8708 5652
rect 9508 5624 9536 5655
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 8680 5596 9536 5624
rect 7577 5587 7635 5593
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 3786 5556 3792 5568
rect 2455 5528 3792 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6914 5556 6920 5568
rect 5776 5528 6920 5556
rect 5776 5516 5782 5528
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7392 5556 7420 5587
rect 8021 5559 8079 5565
rect 8021 5556 8033 5559
rect 7392 5528 8033 5556
rect 8021 5525 8033 5528
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8386 5556 8392 5568
rect 8343 5528 8392 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 9364 5528 9413 5556
rect 9364 5516 9370 5528
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9769 5559 9827 5565
rect 9769 5556 9781 5559
rect 9548 5528 9781 5556
rect 9548 5516 9554 5528
rect 9769 5525 9781 5528
rect 9815 5525 9827 5559
rect 9769 5519 9827 5525
rect 1104 5466 10856 5488
rect 1104 5414 2829 5466
rect 2881 5414 2893 5466
rect 2945 5414 2957 5466
rect 3009 5414 3021 5466
rect 3073 5414 3085 5466
rect 3137 5414 5267 5466
rect 5319 5414 5331 5466
rect 5383 5414 5395 5466
rect 5447 5414 5459 5466
rect 5511 5414 5523 5466
rect 5575 5414 7705 5466
rect 7757 5414 7769 5466
rect 7821 5414 7833 5466
rect 7885 5414 7897 5466
rect 7949 5414 7961 5466
rect 8013 5414 10143 5466
rect 10195 5414 10207 5466
rect 10259 5414 10271 5466
rect 10323 5414 10335 5466
rect 10387 5414 10399 5466
rect 10451 5414 10856 5466
rect 1104 5392 10856 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 3510 5352 3516 5364
rect 2924 5324 3516 5352
rect 2924 5312 2930 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 5261 5355 5319 5361
rect 4264 5324 5028 5352
rect 2317 5287 2375 5293
rect 2317 5284 2329 5287
rect 1688 5256 2329 5284
rect 1688 5228 1716 5256
rect 2317 5253 2329 5256
rect 2363 5284 2375 5287
rect 2363 5256 3280 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1544 5188 1593 5216
rect 1544 5176 1550 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1670 5176 1676 5228
rect 1728 5176 1734 5228
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1780 5188 1869 5216
rect 1780 5148 1808 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 2004 5188 2145 5216
rect 2004 5176 2010 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2222 5176 2228 5228
rect 2280 5176 2286 5228
rect 2498 5176 2504 5228
rect 2556 5176 2562 5228
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5216 2651 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2639 5188 2697 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 3252 5225 3280 5256
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3970 5216 3976 5228
rect 3283 5188 3976 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 2976 5148 3004 5179
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 4172 5160 4200 5312
rect 1596 5120 1808 5148
rect 1872 5120 3004 5148
rect 1596 5092 1624 5120
rect 1578 5040 1584 5092
rect 1636 5040 1642 5092
rect 1872 5089 1900 5120
rect 4154 5108 4160 5160
rect 4212 5108 4218 5160
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5049 1915 5083
rect 1857 5043 1915 5049
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 4264 5080 4292 5324
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5253 4491 5287
rect 4433 5247 4491 5253
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4448 5216 4476 5247
rect 4522 5244 4528 5296
rect 4580 5284 4586 5296
rect 4633 5287 4691 5293
rect 4633 5284 4645 5287
rect 4580 5256 4645 5284
rect 4580 5244 4586 5256
rect 4633 5253 4645 5256
rect 4679 5253 4691 5287
rect 4633 5247 4691 5253
rect 4396 5188 4476 5216
rect 4893 5219 4951 5225
rect 4396 5176 4402 5188
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 5000 5216 5028 5324
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5307 5324 5672 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5644 5293 5672 5324
rect 6546 5312 6552 5364
rect 6604 5312 6610 5364
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5321 9091 5355
rect 9033 5315 9091 5321
rect 5629 5287 5687 5293
rect 5629 5253 5641 5287
rect 5675 5253 5687 5287
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 5629 5247 5687 5253
rect 5736 5256 6377 5284
rect 5736 5216 5764 5256
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6365 5247 6423 5253
rect 5000 5188 5764 5216
rect 5813 5219 5871 5225
rect 4893 5179 4951 5185
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 4908 5148 4936 5179
rect 4356 5120 4936 5148
rect 4985 5151 5043 5157
rect 4356 5089 4384 5120
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 5828 5148 5856 5179
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 5994 5176 6000 5228
rect 6052 5225 6058 5228
rect 6052 5219 6091 5225
rect 6079 5216 6091 5219
rect 6454 5216 6460 5228
rect 6079 5188 6460 5216
rect 6079 5185 6091 5188
rect 6052 5179 6091 5185
rect 6052 5176 6058 5179
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 9048 5216 9076 5315
rect 6687 5188 9076 5216
rect 9401 5219 9459 5225
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9490 5216 9496 5228
rect 9447 5188 9496 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 5828 5120 6408 5148
rect 4985 5111 5043 5117
rect 1995 5052 4292 5080
rect 4341 5083 4399 5089
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 4341 5049 4353 5083
rect 4387 5049 4399 5083
rect 4341 5043 4399 5049
rect 4801 5083 4859 5089
rect 4801 5049 4813 5083
rect 4847 5080 4859 5083
rect 5000 5080 5028 5111
rect 6380 5089 6408 5120
rect 9306 5108 9312 5160
rect 9364 5108 9370 5160
rect 4847 5052 5028 5080
rect 6365 5083 6423 5089
rect 4847 5049 4859 5052
rect 4801 5043 4859 5049
rect 6365 5049 6377 5083
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 2280 4984 3157 5012
rect 2280 4972 2286 4984
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4430 5012 4436 5024
rect 4212 4984 4436 5012
rect 4212 4972 4218 4984
rect 4430 4972 4436 4984
rect 4488 5012 4494 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4488 4984 4629 5012
rect 4488 4972 4494 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 5074 4972 5080 5024
rect 5132 4972 5138 5024
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 10244 5012 10272 5179
rect 5675 4984 10272 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 1854 4808 1860 4820
rect 1627 4780 1860 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 4338 4808 4344 4820
rect 3559 4780 4344 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5074 4768 5080 4820
rect 5132 4768 5138 4820
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 5902 4740 5908 4752
rect 4028 4712 5908 4740
rect 4028 4700 4034 4712
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 4433 4675 4491 4681
rect 3436 4644 4292 4672
rect 3436 4616 3464 4644
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 4264 4604 4292 4644
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 5166 4672 5172 4684
rect 4479 4644 5172 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5224 4644 5365 4672
rect 5224 4632 5230 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 3651 4576 4200 4604
rect 4264 4576 4537 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 3786 4496 3792 4548
rect 3844 4496 3850 4548
rect 3970 4496 3976 4548
rect 4028 4496 4034 4548
rect 4172 4545 4200 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 5276 4536 5304 4567
rect 4203 4508 5304 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 2130 4468 2136 4480
rect 1636 4440 2136 4468
rect 1636 4428 1642 4440
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 4798 4468 4804 4480
rect 3936 4440 4804 4468
rect 3936 4428 3942 4440
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 4890 4428 4896 4480
rect 4948 4428 4954 4480
rect 1104 4378 10856 4400
rect 1104 4326 2829 4378
rect 2881 4326 2893 4378
rect 2945 4326 2957 4378
rect 3009 4326 3021 4378
rect 3073 4326 3085 4378
rect 3137 4326 5267 4378
rect 5319 4326 5331 4378
rect 5383 4326 5395 4378
rect 5447 4326 5459 4378
rect 5511 4326 5523 4378
rect 5575 4326 7705 4378
rect 7757 4326 7769 4378
rect 7821 4326 7833 4378
rect 7885 4326 7897 4378
rect 7949 4326 7961 4378
rect 8013 4326 10143 4378
rect 10195 4326 10207 4378
rect 10259 4326 10271 4378
rect 10323 4326 10335 4378
rect 10387 4326 10399 4378
rect 10451 4326 10856 4378
rect 1104 4304 10856 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1452 4236 2452 4264
rect 1452 4224 1458 4236
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1780 4137 1808 4236
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 2424 4205 2452 4236
rect 2498 4224 2504 4276
rect 2556 4264 2562 4276
rect 2556 4236 2820 4264
rect 2556 4224 2562 4236
rect 2409 4199 2467 4205
rect 2004 4168 2360 4196
rect 2004 4156 2010 4168
rect 2332 4140 2360 4168
rect 2409 4165 2421 4199
rect 2455 4165 2467 4199
rect 2409 4159 2467 4165
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1872 4060 1900 4091
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2314 4088 2320 4140
rect 2372 4088 2378 4140
rect 2498 4088 2504 4140
rect 2556 4088 2562 4140
rect 2792 4137 2820 4236
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3476 4236 3801 4264
rect 3476 4224 3482 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 3789 4227 3847 4233
rect 3510 4196 3516 4208
rect 3068 4168 3516 4196
rect 3068 4137 3096 4168
rect 3510 4156 3516 4168
rect 3568 4156 3574 4208
rect 3804 4196 3832 4227
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5534 4264 5540 4276
rect 4856 4236 5540 4264
rect 4856 4224 4862 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 3804 4168 4568 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 3786 4128 3792 4140
rect 3743 4100 3792 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 2516 4060 2544 4088
rect 1872 4032 2544 4060
rect 2700 4060 2728 4091
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2700 4032 2881 4060
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 3160 3992 3188 4091
rect 3436 4060 3464 4091
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 3970 4128 3976 4140
rect 3927 4100 3976 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 4540 4137 4568 4168
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5132 4168 5580 4196
rect 5132 4156 5138 4168
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 3436 4032 3924 4060
rect 3896 4004 3924 4032
rect 4430 4020 4436 4072
rect 4488 4060 4494 4072
rect 4816 4060 4844 4091
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5552 4137 5580 4168
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 7650 4196 7656 4208
rect 6604 4168 7656 4196
rect 6604 4156 6610 4168
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 7760 4168 8248 4196
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 4948 4100 5273 4128
rect 4948 4088 4954 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 4488 4032 4844 4060
rect 4488 4020 4494 4032
rect 2087 3964 3188 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 3878 3952 3884 4004
rect 3936 3952 3942 4004
rect 1578 3884 1584 3936
rect 1636 3884 1642 3936
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 3234 3924 3240 3936
rect 2179 3896 3240 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 4816 3924 4844 4032
rect 5166 4020 5172 4072
rect 5224 4020 5230 4072
rect 5368 4060 5396 4091
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6638 4128 6644 4140
rect 6328 4100 6644 4128
rect 6328 4088 6334 4100
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6788 4100 6837 4128
rect 6788 4088 6794 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7760 4128 7788 4168
rect 7616 4100 7788 4128
rect 7837 4131 7895 4137
rect 7616 4088 7622 4100
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8110 4128 8116 4140
rect 8067 4100 8116 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 5276 4032 5396 4060
rect 5074 3952 5080 4004
rect 5132 3952 5138 4004
rect 5276 3924 5304 4032
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6420 4032 6561 4060
rect 6420 4020 6426 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 7852 4060 7880 4091
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8220 4128 8248 4168
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8220 4100 8309 4128
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8386 4060 8392 4072
rect 7852 4032 8392 4060
rect 6549 4023 6607 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 4816 3896 5304 3924
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5500 3896 5733 3924
rect 5500 3884 5506 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 7009 3927 7067 3933
rect 7009 3893 7021 3927
rect 7055 3924 7067 3927
rect 7374 3924 7380 3936
rect 7055 3896 7380 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7708 3896 7849 3924
rect 7708 3884 7714 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 8110 3884 8116 3936
rect 8168 3884 8174 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 4430 3680 4436 3732
rect 4488 3680 4494 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 4939 3692 5733 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 4706 3652 4712 3664
rect 1636 3624 4712 3652
rect 1636 3612 1642 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 5074 3652 5080 3664
rect 4847 3624 5080 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 5074 3612 5080 3624
rect 5132 3652 5138 3664
rect 8941 3655 8999 3661
rect 5132 3624 5304 3652
rect 5132 3612 5138 3624
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 1762 3584 1768 3596
rect 1719 3556 1768 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2038 3544 2044 3596
rect 2096 3584 2102 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 2096 3556 2145 3584
rect 2096 3544 2102 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 4985 3587 5043 3593
rect 4985 3553 4997 3587
rect 5031 3584 5043 3587
rect 5166 3584 5172 3596
rect 5031 3556 5172 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1452 3488 2237 3516
rect 1452 3476 1458 3488
rect 2225 3485 2237 3488
rect 2271 3516 2283 3519
rect 3326 3516 3332 3528
rect 2271 3488 3332 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3660 3488 4353 3516
rect 3660 3476 3666 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 5276 3525 5304 3624
rect 5368 3624 8524 3652
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 842 3408 848 3460
rect 900 3448 906 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 900 3420 1501 3448
rect 900 3408 906 3420
rect 1489 3417 1501 3420
rect 1535 3417 1547 3451
rect 1489 3411 1547 3417
rect 5077 3451 5135 3457
rect 5077 3417 5089 3451
rect 5123 3448 5135 3451
rect 5368 3448 5396 3624
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6380 3556 6837 3584
rect 6380 3528 6408 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 7006 3544 7012 3596
rect 7064 3544 7070 3596
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 8205 3587 8263 3593
rect 7239 3556 7328 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 6362 3476 6368 3528
rect 6420 3476 6426 3528
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 6914 3476 6920 3528
rect 6972 3476 6978 3528
rect 7300 3525 7328 3556
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8386 3584 8392 3596
rect 8251 3556 8392 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8496 3516 8524 3624
rect 8941 3621 8953 3655
rect 8987 3652 8999 3655
rect 8987 3624 10272 3652
rect 8987 3621 8999 3624
rect 8941 3615 8999 3621
rect 9398 3584 9404 3596
rect 9329 3556 9404 3584
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8496 3488 9137 3516
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9329 3503 9357 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 10244 3525 10272 3624
rect 10229 3519 10287 3525
rect 9125 3479 9183 3485
rect 9314 3497 9372 3503
rect 9314 3463 9326 3497
rect 9360 3463 9372 3497
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 5123 3420 5396 3448
rect 5123 3417 5135 3420
rect 5077 3411 5135 3417
rect 5534 3408 5540 3460
rect 5592 3408 5598 3460
rect 5644 3420 8156 3448
rect 2590 3340 2596 3392
rect 2648 3340 2654 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 5644 3380 5672 3420
rect 8128 3392 8156 3420
rect 8938 3408 8944 3460
rect 8996 3408 9002 3460
rect 9214 3408 9220 3460
rect 9272 3408 9278 3460
rect 9314 3457 9372 3463
rect 3292 3352 5672 3380
rect 3292 3340 3298 3352
rect 5718 3340 5724 3392
rect 5776 3389 5782 3392
rect 5776 3383 5795 3389
rect 5783 3349 5795 3383
rect 5776 3343 5795 3349
rect 5776 3340 5782 3343
rect 5902 3340 5908 3392
rect 5960 3340 5966 3392
rect 5994 3340 6000 3392
rect 6052 3340 6058 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 6880 3352 7849 3380
rect 6880 3340 6886 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 7837 3343 7895 3349
rect 8110 3340 8116 3392
rect 8168 3340 8174 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8481 3383 8539 3389
rect 8481 3380 8493 3383
rect 8444 3352 8493 3380
rect 8444 3340 8450 3352
rect 8481 3349 8493 3352
rect 8527 3349 8539 3383
rect 8481 3343 8539 3349
rect 10413 3383 10471 3389
rect 10413 3349 10425 3383
rect 10459 3380 10471 3383
rect 10502 3380 10508 3392
rect 10459 3352 10508 3380
rect 10459 3349 10471 3352
rect 10413 3343 10471 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 1104 3290 10856 3312
rect 1104 3238 2829 3290
rect 2881 3238 2893 3290
rect 2945 3238 2957 3290
rect 3009 3238 3021 3290
rect 3073 3238 3085 3290
rect 3137 3238 5267 3290
rect 5319 3238 5331 3290
rect 5383 3238 5395 3290
rect 5447 3238 5459 3290
rect 5511 3238 5523 3290
rect 5575 3238 7705 3290
rect 7757 3238 7769 3290
rect 7821 3238 7833 3290
rect 7885 3238 7897 3290
rect 7949 3238 7961 3290
rect 8013 3238 10143 3290
rect 10195 3238 10207 3290
rect 10259 3238 10271 3290
rect 10323 3238 10335 3290
rect 10387 3238 10399 3290
rect 10451 3238 10856 3290
rect 1104 3216 10856 3238
rect 1946 3136 1952 3188
rect 2004 3136 2010 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4706 3176 4712 3188
rect 4203 3148 4712 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4706 3136 4712 3148
rect 4764 3176 4770 3188
rect 5258 3176 5264 3188
rect 4764 3148 5264 3176
rect 4764 3136 4770 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5718 3176 5724 3188
rect 5583 3148 5724 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5994 3176 6000 3188
rect 5828 3148 6000 3176
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 2498 3108 2504 3120
rect 1719 3080 2504 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 2498 3068 2504 3080
rect 2556 3108 2562 3120
rect 5828 3108 5856 3148
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 6788 3148 7205 3176
rect 6788 3136 6794 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 8211 3179 8269 3185
rect 8211 3145 8223 3179
rect 8257 3176 8269 3179
rect 8938 3176 8944 3188
rect 8257 3148 8944 3176
rect 8257 3145 8269 3148
rect 8211 3139 8269 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 2556 3080 3924 3108
rect 2556 3068 2562 3080
rect 1486 3000 1492 3052
rect 1544 3000 1550 3052
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 3252 3049 3280 3080
rect 3896 3052 3924 3080
rect 4540 3080 5856 3108
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 3145 2975 3203 2981
rect 3145 2972 3157 2975
rect 2648 2944 3157 2972
rect 2648 2932 2654 2944
rect 3145 2941 3157 2944
rect 3191 2972 3203 2975
rect 3712 2972 3740 3003
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 4540 3049 4568 3080
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 5960 3080 6776 3108
rect 5960 3068 5966 3080
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 5166 3040 5172 3052
rect 4525 3003 4583 3009
rect 4908 3012 5172 3040
rect 3191 2944 3740 2972
rect 3789 2975 3847 2981
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 4080 2972 4108 3003
rect 3835 2944 4108 2972
rect 4617 2975 4675 2981
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4798 2972 4804 2984
rect 4663 2944 4804 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 4908 2981 4936 3012
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 6748 3049 6776 3080
rect 6932 3080 7481 3108
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 6932 3049 6960 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 8110 3068 8116 3120
rect 8168 3068 8174 3120
rect 9398 3108 9404 3120
rect 8220 3080 9404 3108
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 5132 2944 5212 2972
rect 5132 2932 5138 2944
rect 3602 2864 3608 2916
rect 3660 2864 3666 2916
rect 5184 2836 5212 2944
rect 5258 2932 5264 2984
rect 5316 2932 5322 2984
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2972 6515 2975
rect 7006 2972 7012 2984
rect 6503 2944 7012 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 7116 2904 7144 3003
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7742 3040 7748 3052
rect 7607 3012 7748 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7392 2972 7420 3003
rect 7742 3000 7748 3012
rect 7800 3040 7806 3052
rect 8220 3040 8248 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 7800 3012 8248 3040
rect 8297 3043 8355 3049
rect 7800 3000 7806 3012
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 6052 2876 7144 2904
rect 7300 2944 7420 2972
rect 6052 2864 6058 2876
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 5184 2808 5273 2836
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5261 2799 5319 2805
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 7300 2836 7328 2944
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8312 2972 8340 3003
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 7708 2944 8340 2972
rect 7708 2932 7714 2944
rect 6420 2808 7328 2836
rect 6420 2796 6426 2808
rect 7374 2796 7380 2848
rect 7432 2836 7438 2848
rect 10226 2836 10232 2848
rect 7432 2808 10232 2836
rect 7432 2796 7438 2808
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 1670 2456 1676 2508
rect 1728 2456 1734 2508
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 10226 2388 10232 2440
rect 10284 2388 10290 2440
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 9640 2264 10425 2292
rect 9640 2252 9646 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 1104 2202 10856 2224
rect 1104 2150 2829 2202
rect 2881 2150 2893 2202
rect 2945 2150 2957 2202
rect 3009 2150 3021 2202
rect 3073 2150 3085 2202
rect 3137 2150 5267 2202
rect 5319 2150 5331 2202
rect 5383 2150 5395 2202
rect 5447 2150 5459 2202
rect 5511 2150 5523 2202
rect 5575 2150 7705 2202
rect 7757 2150 7769 2202
rect 7821 2150 7833 2202
rect 7885 2150 7897 2202
rect 7949 2150 7961 2202
rect 8013 2150 10143 2202
rect 10195 2150 10207 2202
rect 10259 2150 10271 2202
rect 10323 2150 10335 2202
rect 10387 2150 10399 2202
rect 10451 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 2169 13574 2221 13626
rect 2233 13574 2285 13626
rect 2297 13574 2349 13626
rect 2361 13574 2413 13626
rect 2425 13574 2477 13626
rect 4607 13574 4659 13626
rect 4671 13574 4723 13626
rect 4735 13574 4787 13626
rect 4799 13574 4851 13626
rect 4863 13574 4915 13626
rect 7045 13574 7097 13626
rect 7109 13574 7161 13626
rect 7173 13574 7225 13626
rect 7237 13574 7289 13626
rect 7301 13574 7353 13626
rect 9483 13574 9535 13626
rect 9547 13574 9599 13626
rect 9611 13574 9663 13626
rect 9675 13574 9727 13626
rect 9739 13574 9791 13626
rect 10416 13515 10468 13524
rect 10416 13481 10425 13515
rect 10425 13481 10459 13515
rect 10459 13481 10468 13515
rect 10416 13472 10468 13481
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2228 13268 2280 13320
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 3608 13311 3660 13320
rect 3608 13277 3617 13311
rect 3617 13277 3651 13311
rect 3651 13277 3660 13311
rect 3608 13268 3660 13277
rect 8576 13268 8628 13320
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 3516 13200 3568 13252
rect 1400 13132 1452 13184
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 3332 13132 3384 13184
rect 2829 13030 2881 13082
rect 2893 13030 2945 13082
rect 2957 13030 3009 13082
rect 3021 13030 3073 13082
rect 3085 13030 3137 13082
rect 5267 13030 5319 13082
rect 5331 13030 5383 13082
rect 5395 13030 5447 13082
rect 5459 13030 5511 13082
rect 5523 13030 5575 13082
rect 7705 13030 7757 13082
rect 7769 13030 7821 13082
rect 7833 13030 7885 13082
rect 7897 13030 7949 13082
rect 7961 13030 8013 13082
rect 10143 13030 10195 13082
rect 10207 13030 10259 13082
rect 10271 13030 10323 13082
rect 10335 13030 10387 13082
rect 10399 13030 10451 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 2596 12928 2648 12980
rect 4988 12928 5040 12980
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 3240 12860 3292 12912
rect 2504 12724 2556 12776
rect 2872 12792 2924 12844
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 5172 12724 5224 12776
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 6276 12724 6328 12776
rect 7932 12792 7984 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 7380 12724 7432 12776
rect 5540 12656 5592 12708
rect 8576 12656 8628 12708
rect 2044 12588 2096 12597
rect 4528 12588 4580 12640
rect 6828 12588 6880 12640
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 7472 12588 7524 12640
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 2169 12486 2221 12538
rect 2233 12486 2285 12538
rect 2297 12486 2349 12538
rect 2361 12486 2413 12538
rect 2425 12486 2477 12538
rect 4607 12486 4659 12538
rect 4671 12486 4723 12538
rect 4735 12486 4787 12538
rect 4799 12486 4851 12538
rect 4863 12486 4915 12538
rect 7045 12486 7097 12538
rect 7109 12486 7161 12538
rect 7173 12486 7225 12538
rect 7237 12486 7289 12538
rect 7301 12486 7353 12538
rect 9483 12486 9535 12538
rect 9547 12486 9599 12538
rect 9611 12486 9663 12538
rect 9675 12486 9727 12538
rect 9739 12486 9791 12538
rect 1952 12384 2004 12436
rect 1676 12316 1728 12368
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 2688 12316 2740 12368
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2688 12180 2740 12232
rect 3332 12384 3384 12436
rect 3976 12316 4028 12368
rect 4436 12316 4488 12368
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 3516 12248 3568 12300
rect 1492 12112 1544 12164
rect 1952 12112 2004 12164
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3424 12180 3476 12232
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 4160 12180 4212 12232
rect 3608 12112 3660 12164
rect 4712 12316 4764 12368
rect 4896 12248 4948 12300
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5908 12316 5960 12368
rect 6092 12359 6144 12368
rect 6092 12325 6101 12359
rect 6101 12325 6135 12359
rect 6135 12325 6144 12359
rect 6092 12316 6144 12325
rect 5816 12248 5868 12300
rect 4160 12044 4212 12096
rect 4804 12044 4856 12096
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 6920 12316 6972 12368
rect 7012 12316 7064 12368
rect 7748 12316 7800 12368
rect 7932 12316 7984 12368
rect 6552 12180 6604 12232
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7564 12180 7616 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 5632 12044 5684 12096
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 6920 12044 6972 12096
rect 7288 12155 7340 12164
rect 7288 12121 7323 12155
rect 7323 12121 7340 12155
rect 7288 12112 7340 12121
rect 7932 12155 7984 12164
rect 7932 12121 7941 12155
rect 7941 12121 7975 12155
rect 7975 12121 7984 12155
rect 7932 12112 7984 12121
rect 8208 12044 8260 12096
rect 9312 12044 9364 12096
rect 2829 11942 2881 11994
rect 2893 11942 2945 11994
rect 2957 11942 3009 11994
rect 3021 11942 3073 11994
rect 3085 11942 3137 11994
rect 5267 11942 5319 11994
rect 5331 11942 5383 11994
rect 5395 11942 5447 11994
rect 5459 11942 5511 11994
rect 5523 11942 5575 11994
rect 7705 11942 7757 11994
rect 7769 11942 7821 11994
rect 7833 11942 7885 11994
rect 7897 11942 7949 11994
rect 7961 11942 8013 11994
rect 10143 11942 10195 11994
rect 10207 11942 10259 11994
rect 10271 11942 10323 11994
rect 10335 11942 10387 11994
rect 10399 11942 10451 11994
rect 2504 11840 2556 11892
rect 2688 11840 2740 11892
rect 1860 11772 1912 11824
rect 2964 11772 3016 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 2044 11704 2096 11756
rect 3240 11704 3292 11756
rect 3884 11840 3936 11892
rect 4988 11883 5040 11892
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5172 11840 5224 11892
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 4436 11772 4488 11824
rect 4712 11772 4764 11824
rect 3976 11636 4028 11688
rect 2872 11568 2924 11620
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 4344 11704 4396 11756
rect 4988 11704 5040 11756
rect 6000 11772 6052 11824
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 7472 11840 7524 11892
rect 7748 11840 7800 11892
rect 6920 11704 6972 11756
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8300 11772 8352 11824
rect 10232 11772 10284 11824
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 3148 11500 3200 11552
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 4160 11568 4212 11620
rect 4252 11568 4304 11620
rect 5264 11568 5316 11620
rect 4436 11500 4488 11552
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 4804 11500 4856 11552
rect 5172 11500 5224 11552
rect 6184 11568 6236 11620
rect 8392 11636 8444 11688
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 6644 11500 6696 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8116 11500 8168 11552
rect 9864 11500 9916 11552
rect 2169 11398 2221 11450
rect 2233 11398 2285 11450
rect 2297 11398 2349 11450
rect 2361 11398 2413 11450
rect 2425 11398 2477 11450
rect 4607 11398 4659 11450
rect 4671 11398 4723 11450
rect 4735 11398 4787 11450
rect 4799 11398 4851 11450
rect 4863 11398 4915 11450
rect 7045 11398 7097 11450
rect 7109 11398 7161 11450
rect 7173 11398 7225 11450
rect 7237 11398 7289 11450
rect 7301 11398 7353 11450
rect 9483 11398 9535 11450
rect 9547 11398 9599 11450
rect 9611 11398 9663 11450
rect 9675 11398 9727 11450
rect 9739 11398 9791 11450
rect 2596 11296 2648 11348
rect 3424 11296 3476 11348
rect 4160 11296 4212 11348
rect 4988 11296 5040 11348
rect 6368 11296 6420 11348
rect 7472 11296 7524 11348
rect 8024 11296 8076 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 2320 11228 2372 11280
rect 3240 11228 3292 11280
rect 3792 11228 3844 11280
rect 4344 11228 4396 11280
rect 4436 11228 4488 11280
rect 4804 11228 4856 11280
rect 848 11092 900 11144
rect 1584 11092 1636 11144
rect 1860 11092 1912 11144
rect 2596 11092 2648 11144
rect 3148 11092 3200 11144
rect 3240 11092 3292 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4252 11160 4304 11212
rect 4528 11160 4580 11212
rect 4160 11092 4212 11144
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 2044 11024 2096 11076
rect 2320 11024 2372 11076
rect 2872 11024 2924 11076
rect 3516 11024 3568 11076
rect 4528 11024 4580 11076
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 6920 11160 6972 11212
rect 6552 11092 6604 11144
rect 7932 11228 7984 11280
rect 8208 11271 8260 11280
rect 8208 11237 8217 11271
rect 8217 11237 8251 11271
rect 8251 11237 8260 11271
rect 8208 11228 8260 11237
rect 9772 11296 9824 11348
rect 10048 11228 10100 11280
rect 10232 11271 10284 11280
rect 10232 11237 10241 11271
rect 10241 11237 10275 11271
rect 10275 11237 10284 11271
rect 10232 11228 10284 11237
rect 10508 11228 10560 11280
rect 9128 11160 9180 11212
rect 9772 11160 9824 11212
rect 2964 10956 3016 11008
rect 4068 10956 4120 11008
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 7748 11024 7800 11076
rect 7564 10956 7616 11008
rect 8024 11024 8076 11076
rect 9864 11067 9916 11076
rect 9864 11033 9873 11067
rect 9873 11033 9907 11067
rect 9907 11033 9916 11067
rect 9864 11024 9916 11033
rect 9036 10956 9088 11008
rect 2829 10854 2881 10906
rect 2893 10854 2945 10906
rect 2957 10854 3009 10906
rect 3021 10854 3073 10906
rect 3085 10854 3137 10906
rect 5267 10854 5319 10906
rect 5331 10854 5383 10906
rect 5395 10854 5447 10906
rect 5459 10854 5511 10906
rect 5523 10854 5575 10906
rect 7705 10854 7757 10906
rect 7769 10854 7821 10906
rect 7833 10854 7885 10906
rect 7897 10854 7949 10906
rect 7961 10854 8013 10906
rect 10143 10854 10195 10906
rect 10207 10854 10259 10906
rect 10271 10854 10323 10906
rect 10335 10854 10387 10906
rect 10399 10854 10451 10906
rect 4620 10752 4672 10804
rect 848 10616 900 10668
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 5264 10752 5316 10804
rect 5724 10752 5776 10804
rect 6000 10752 6052 10804
rect 6276 10752 6328 10804
rect 9036 10752 9088 10804
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 4160 10548 4212 10600
rect 1952 10480 2004 10532
rect 4896 10480 4948 10532
rect 1860 10455 1912 10464
rect 1860 10421 1869 10455
rect 1869 10421 1903 10455
rect 1903 10421 1912 10455
rect 1860 10412 1912 10421
rect 4344 10455 4396 10464
rect 4344 10421 4353 10455
rect 4353 10421 4387 10455
rect 4387 10421 4396 10455
rect 4344 10412 4396 10421
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 7380 10684 7432 10736
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6000 10548 6052 10557
rect 5448 10480 5500 10532
rect 6920 10616 6972 10668
rect 7472 10616 7524 10668
rect 7564 10616 7616 10668
rect 6184 10548 6236 10600
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 10048 10616 10100 10668
rect 8208 10480 8260 10532
rect 6000 10412 6052 10464
rect 8944 10412 8996 10464
rect 2169 10310 2221 10362
rect 2233 10310 2285 10362
rect 2297 10310 2349 10362
rect 2361 10310 2413 10362
rect 2425 10310 2477 10362
rect 4607 10310 4659 10362
rect 4671 10310 4723 10362
rect 4735 10310 4787 10362
rect 4799 10310 4851 10362
rect 4863 10310 4915 10362
rect 7045 10310 7097 10362
rect 7109 10310 7161 10362
rect 7173 10310 7225 10362
rect 7237 10310 7289 10362
rect 7301 10310 7353 10362
rect 9483 10310 9535 10362
rect 9547 10310 9599 10362
rect 9611 10310 9663 10362
rect 9675 10310 9727 10362
rect 9739 10310 9791 10362
rect 2964 10208 3016 10260
rect 3976 10208 4028 10260
rect 5172 10208 5224 10260
rect 5816 10208 5868 10260
rect 1860 10140 1912 10192
rect 6552 10140 6604 10192
rect 8760 10140 8812 10192
rect 3884 10072 3936 10124
rect 3976 10072 4028 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 1492 9979 1544 9988
rect 1492 9945 1501 9979
rect 1501 9945 1535 9979
rect 1535 9945 1544 9979
rect 1492 9936 1544 9945
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 2044 9936 2096 9988
rect 2688 9936 2740 9988
rect 3332 10004 3384 10056
rect 6000 10072 6052 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 6000 9936 6052 9988
rect 1860 9868 1912 9920
rect 2872 9868 2924 9920
rect 3516 9868 3568 9920
rect 6644 9868 6696 9920
rect 9680 9868 9732 9920
rect 2829 9766 2881 9818
rect 2893 9766 2945 9818
rect 2957 9766 3009 9818
rect 3021 9766 3073 9818
rect 3085 9766 3137 9818
rect 5267 9766 5319 9818
rect 5331 9766 5383 9818
rect 5395 9766 5447 9818
rect 5459 9766 5511 9818
rect 5523 9766 5575 9818
rect 7705 9766 7757 9818
rect 7769 9766 7821 9818
rect 7833 9766 7885 9818
rect 7897 9766 7949 9818
rect 7961 9766 8013 9818
rect 10143 9766 10195 9818
rect 10207 9766 10259 9818
rect 10271 9766 10323 9818
rect 10335 9766 10387 9818
rect 10399 9766 10451 9818
rect 1768 9664 1820 9716
rect 2596 9664 2648 9716
rect 2780 9596 2832 9648
rect 3976 9664 4028 9716
rect 4160 9707 4212 9716
rect 4160 9673 4169 9707
rect 4169 9673 4203 9707
rect 4203 9673 4212 9707
rect 4160 9664 4212 9673
rect 1860 9528 1912 9580
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 1768 9460 1820 9512
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 3240 9528 3292 9580
rect 3148 9460 3200 9512
rect 4068 9596 4120 9648
rect 6552 9639 6604 9648
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 6184 9528 6236 9580
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 3976 9460 4028 9512
rect 4988 9460 5040 9512
rect 6092 9460 6144 9512
rect 8116 9596 8168 9648
rect 6828 9528 6880 9580
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 4068 9392 4120 9444
rect 5356 9392 5408 9444
rect 6920 9460 6972 9512
rect 8024 9460 8076 9512
rect 8944 9460 8996 9512
rect 8300 9392 8352 9444
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 3148 9324 3200 9376
rect 3240 9324 3292 9376
rect 6276 9324 6328 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 9312 9324 9364 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 1952 9120 2004 9172
rect 3240 9120 3292 9172
rect 3884 9120 3936 9172
rect 3516 9052 3568 9104
rect 848 8916 900 8968
rect 1492 8916 1544 8968
rect 2504 8916 2556 8968
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3792 8984 3844 9036
rect 5540 9052 5592 9104
rect 6092 9052 6144 9104
rect 7012 9120 7064 9172
rect 8760 9120 8812 9172
rect 6736 9052 6788 9104
rect 6920 9095 6972 9104
rect 6920 9061 6929 9095
rect 6929 9061 6963 9095
rect 6963 9061 6972 9095
rect 6920 9052 6972 9061
rect 5724 8959 5776 8968
rect 1860 8848 1912 8900
rect 5724 8925 5738 8959
rect 5738 8925 5772 8959
rect 5772 8925 5776 8959
rect 5724 8916 5776 8925
rect 5356 8891 5408 8900
rect 5356 8857 5365 8891
rect 5365 8857 5399 8891
rect 5399 8857 5408 8891
rect 5356 8848 5408 8857
rect 5540 8891 5592 8900
rect 5540 8857 5549 8891
rect 5549 8857 5583 8891
rect 5583 8857 5592 8891
rect 5540 8848 5592 8857
rect 2044 8780 2096 8832
rect 4068 8780 4120 8832
rect 4344 8780 4396 8832
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6092 8891 6144 8900
rect 6092 8857 6101 8891
rect 6101 8857 6135 8891
rect 6135 8857 6144 8891
rect 6092 8848 6144 8857
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 6644 8916 6696 8968
rect 7380 8916 7432 8968
rect 7104 8848 7156 8900
rect 7288 8848 7340 8900
rect 6552 8780 6604 8832
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 7196 8780 7248 8832
rect 7564 8848 7616 8900
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 8300 8916 8352 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 10048 8984 10100 9036
rect 8116 8823 8168 8832
rect 8116 8789 8125 8823
rect 8125 8789 8159 8823
rect 8159 8789 8168 8823
rect 8116 8780 8168 8789
rect 8208 8780 8260 8832
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10048 8848 10100 8900
rect 9864 8780 9916 8832
rect 2829 8678 2881 8730
rect 2893 8678 2945 8730
rect 2957 8678 3009 8730
rect 3021 8678 3073 8730
rect 3085 8678 3137 8730
rect 5267 8678 5319 8730
rect 5331 8678 5383 8730
rect 5395 8678 5447 8730
rect 5459 8678 5511 8730
rect 5523 8678 5575 8730
rect 7705 8678 7757 8730
rect 7769 8678 7821 8730
rect 7833 8678 7885 8730
rect 7897 8678 7949 8730
rect 7961 8678 8013 8730
rect 10143 8678 10195 8730
rect 10207 8678 10259 8730
rect 10271 8678 10323 8730
rect 10335 8678 10387 8730
rect 10399 8678 10451 8730
rect 7288 8619 7340 8628
rect 7288 8585 7297 8619
rect 7297 8585 7331 8619
rect 7331 8585 7340 8619
rect 7288 8576 7340 8585
rect 7564 8576 7616 8628
rect 8208 8576 8260 8628
rect 3240 8440 3292 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 1768 8372 1820 8424
rect 4620 8440 4672 8492
rect 6460 8551 6512 8560
rect 6460 8517 6469 8551
rect 6469 8517 6503 8551
rect 6503 8517 6512 8551
rect 6460 8508 6512 8517
rect 6644 8551 6696 8560
rect 6644 8517 6653 8551
rect 6653 8517 6687 8551
rect 6687 8517 6696 8551
rect 10876 8576 10928 8628
rect 6644 8508 6696 8517
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6276 8440 6328 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7104 8372 7156 8424
rect 7288 8440 7340 8492
rect 7472 8440 7524 8492
rect 8024 8372 8076 8424
rect 4160 8236 4212 8288
rect 4620 8304 4672 8356
rect 4436 8236 4488 8288
rect 6736 8304 6788 8356
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 5632 8236 5684 8288
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 9864 8440 9916 8492
rect 10048 8440 10100 8492
rect 8392 8236 8444 8245
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 1676 8032 1728 8084
rect 2044 8007 2096 8016
rect 2044 7973 2053 8007
rect 2053 7973 2087 8007
rect 2087 7973 2096 8007
rect 2044 7964 2096 7973
rect 2596 8032 2648 8084
rect 2688 7964 2740 8016
rect 2504 7828 2556 7880
rect 4712 8032 4764 8084
rect 5080 8032 5132 8084
rect 5632 8032 5684 8084
rect 6460 8032 6512 8084
rect 4620 7964 4672 8016
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4528 7828 4580 7880
rect 6000 7896 6052 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 6828 7896 6880 7948
rect 7380 7896 7432 7948
rect 2596 7760 2648 7812
rect 5080 7760 5132 7812
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 3884 7692 3936 7744
rect 7564 7828 7616 7880
rect 7472 7692 7524 7744
rect 2829 7590 2881 7642
rect 2893 7590 2945 7642
rect 2957 7590 3009 7642
rect 3021 7590 3073 7642
rect 3085 7590 3137 7642
rect 5267 7590 5319 7642
rect 5331 7590 5383 7642
rect 5395 7590 5447 7642
rect 5459 7590 5511 7642
rect 5523 7590 5575 7642
rect 7705 7590 7757 7642
rect 7769 7590 7821 7642
rect 7833 7590 7885 7642
rect 7897 7590 7949 7642
rect 7961 7590 8013 7642
rect 10143 7590 10195 7642
rect 10207 7590 10259 7642
rect 10271 7590 10323 7642
rect 10335 7590 10387 7642
rect 10399 7590 10451 7642
rect 1400 7488 1452 7540
rect 1768 7420 1820 7472
rect 848 7352 900 7404
rect 1676 7352 1728 7404
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 4436 7488 4488 7540
rect 4988 7488 5040 7540
rect 2596 7420 2648 7472
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 3240 7284 3292 7336
rect 4160 7352 4212 7404
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 2044 7148 2096 7200
rect 2412 7148 2464 7200
rect 4436 7216 4488 7268
rect 4620 7216 4672 7268
rect 6000 7216 6052 7268
rect 2780 7148 2832 7200
rect 4160 7148 4212 7200
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4712 7148 4764 7200
rect 5080 7148 5132 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 2780 6944 2832 6996
rect 2412 6876 2464 6928
rect 2688 6876 2740 6928
rect 848 6740 900 6792
rect 1584 6740 1636 6792
rect 1768 6740 1820 6792
rect 1952 6715 2004 6724
rect 1952 6681 1961 6715
rect 1961 6681 1995 6715
rect 1995 6681 2004 6715
rect 1952 6672 2004 6681
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 4160 6876 4212 6928
rect 4620 6876 4672 6928
rect 5724 6944 5776 6996
rect 10232 6944 10284 6996
rect 6644 6876 6696 6928
rect 3976 6808 4028 6860
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 3424 6672 3476 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 1676 6604 1728 6656
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 4436 6672 4488 6724
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 5264 6715 5316 6724
rect 5264 6681 5273 6715
rect 5273 6681 5307 6715
rect 5307 6681 5316 6715
rect 5264 6672 5316 6681
rect 5632 6740 5684 6792
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6368 6740 6420 6792
rect 8116 6808 8168 6860
rect 9036 6876 9088 6928
rect 9496 6876 9548 6928
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7564 6740 7616 6792
rect 8392 6740 8444 6792
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9220 6740 9272 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 10048 6740 10100 6792
rect 6736 6672 6788 6724
rect 7472 6604 7524 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 8668 6604 8720 6656
rect 9772 6604 9824 6656
rect 2829 6502 2881 6554
rect 2893 6502 2945 6554
rect 2957 6502 3009 6554
rect 3021 6502 3073 6554
rect 3085 6502 3137 6554
rect 5267 6502 5319 6554
rect 5331 6502 5383 6554
rect 5395 6502 5447 6554
rect 5459 6502 5511 6554
rect 5523 6502 5575 6554
rect 7705 6502 7757 6554
rect 7769 6502 7821 6554
rect 7833 6502 7885 6554
rect 7897 6502 7949 6554
rect 7961 6502 8013 6554
rect 10143 6502 10195 6554
rect 10207 6502 10259 6554
rect 10271 6502 10323 6554
rect 10335 6502 10387 6554
rect 10399 6502 10451 6554
rect 1584 6400 1636 6452
rect 3332 6400 3384 6452
rect 4712 6400 4764 6452
rect 5816 6400 5868 6452
rect 1952 6332 2004 6384
rect 3240 6375 3292 6384
rect 3240 6341 3249 6375
rect 3249 6341 3283 6375
rect 3283 6341 3292 6375
rect 3240 6332 3292 6341
rect 1584 6264 1636 6316
rect 1768 6264 1820 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 4160 6332 4212 6384
rect 4896 6332 4948 6384
rect 6368 6400 6420 6452
rect 7472 6400 7524 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 1952 6196 2004 6248
rect 2228 6196 2280 6248
rect 4068 6196 4120 6248
rect 5632 6196 5684 6248
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 6184 6264 6236 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7840 6332 7892 6384
rect 8116 6264 8168 6316
rect 8944 6264 8996 6316
rect 7380 6196 7432 6248
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 7656 6196 7708 6248
rect 6000 6128 6052 6180
rect 6276 6128 6328 6180
rect 6828 6128 6880 6180
rect 7288 6128 7340 6180
rect 7840 6128 7892 6180
rect 9220 6196 9272 6248
rect 9864 6264 9916 6316
rect 9956 6196 10008 6248
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 2596 6060 2648 6112
rect 4344 6060 4396 6112
rect 7380 6060 7432 6112
rect 8300 6060 8352 6112
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 6828 5856 6880 5908
rect 7380 5856 7432 5908
rect 6000 5788 6052 5840
rect 7748 5831 7800 5840
rect 7748 5797 7757 5831
rect 7757 5797 7791 5831
rect 7791 5797 7800 5831
rect 7748 5788 7800 5797
rect 7932 5788 7984 5840
rect 8208 5788 8260 5840
rect 2504 5720 2556 5772
rect 6092 5720 6144 5772
rect 7472 5720 7524 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1492 5652 1544 5704
rect 2228 5652 2280 5704
rect 4344 5652 4396 5704
rect 6920 5652 6972 5704
rect 6276 5584 6328 5636
rect 8300 5652 8352 5704
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 3792 5516 3844 5568
rect 5724 5516 5776 5568
rect 6920 5516 6972 5568
rect 8392 5516 8444 5568
rect 9312 5516 9364 5568
rect 9496 5516 9548 5568
rect 2829 5414 2881 5466
rect 2893 5414 2945 5466
rect 2957 5414 3009 5466
rect 3021 5414 3073 5466
rect 3085 5414 3137 5466
rect 5267 5414 5319 5466
rect 5331 5414 5383 5466
rect 5395 5414 5447 5466
rect 5459 5414 5511 5466
rect 5523 5414 5575 5466
rect 7705 5414 7757 5466
rect 7769 5414 7821 5466
rect 7833 5414 7885 5466
rect 7897 5414 7949 5466
rect 7961 5414 8013 5466
rect 10143 5414 10195 5466
rect 10207 5414 10259 5466
rect 10271 5414 10323 5466
rect 10335 5414 10387 5466
rect 10399 5414 10451 5466
rect 2872 5312 2924 5364
rect 3516 5312 3568 5364
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 1492 5176 1544 5228
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 1952 5176 2004 5228
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3976 5176 4028 5228
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 1584 5040 1636 5092
rect 4160 5108 4212 5160
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4528 5244 4580 5296
rect 4344 5176 4396 5185
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6000 5219 6052 5228
rect 6000 5185 6045 5219
rect 6045 5185 6052 5219
rect 6000 5176 6052 5185
rect 6460 5176 6512 5228
rect 9496 5176 9548 5228
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 2228 4972 2280 5024
rect 4160 4972 4212 5024
rect 4436 4972 4488 5024
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 5080 4972 5132 4981
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 1860 4768 1912 4820
rect 4344 4768 4396 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 3976 4700 4028 4752
rect 5908 4700 5960 4752
rect 848 4564 900 4616
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 5172 4632 5224 4684
rect 3792 4539 3844 4548
rect 3792 4505 3801 4539
rect 3801 4505 3835 4539
rect 3835 4505 3844 4539
rect 3792 4496 3844 4505
rect 3976 4539 4028 4548
rect 3976 4505 3985 4539
rect 3985 4505 4019 4539
rect 4019 4505 4028 4539
rect 3976 4496 4028 4505
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4804 4564 4856 4616
rect 1584 4428 1636 4480
rect 2136 4428 2188 4480
rect 3884 4428 3936 4480
rect 4804 4428 4856 4480
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 2829 4326 2881 4378
rect 2893 4326 2945 4378
rect 2957 4326 3009 4378
rect 3021 4326 3073 4378
rect 3085 4326 3137 4378
rect 5267 4326 5319 4378
rect 5331 4326 5383 4378
rect 5395 4326 5447 4378
rect 5459 4326 5511 4378
rect 5523 4326 5575 4378
rect 7705 4326 7757 4378
rect 7769 4326 7821 4378
rect 7833 4326 7885 4378
rect 7897 4326 7949 4378
rect 7961 4326 8013 4378
rect 10143 4326 10195 4378
rect 10207 4326 10259 4378
rect 10271 4326 10323 4378
rect 10335 4326 10387 4378
rect 10399 4326 10451 4378
rect 1400 4224 1452 4276
rect 848 4088 900 4140
rect 1952 4156 2004 4208
rect 2504 4224 2556 4276
rect 2136 4088 2188 4140
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 3424 4224 3476 4276
rect 3516 4156 3568 4208
rect 4804 4224 4856 4276
rect 5540 4224 5592 4276
rect 3792 4088 3844 4140
rect 3976 4088 4028 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 5080 4156 5132 4208
rect 4436 4020 4488 4072
rect 4896 4088 4948 4140
rect 6552 4156 6604 4208
rect 7656 4156 7708 4208
rect 3884 3952 3936 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 3240 3884 3292 3936
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 6276 4088 6328 4140
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6736 4088 6788 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 8116 4131 8168 4140
rect 5080 3995 5132 4004
rect 5080 3961 5089 3995
rect 5089 3961 5123 3995
rect 5123 3961 5132 3995
rect 5080 3952 5132 3961
rect 6368 4020 6420 4072
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8392 4020 8444 4072
rect 5448 3884 5500 3936
rect 7380 3884 7432 3936
rect 7656 3884 7708 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 1584 3612 1636 3664
rect 4712 3612 4764 3664
rect 5080 3612 5132 3664
rect 1768 3544 1820 3596
rect 2044 3544 2096 3596
rect 5172 3544 5224 3596
rect 1400 3476 1452 3528
rect 3332 3476 3384 3528
rect 3608 3476 3660 3528
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 848 3408 900 3460
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 8392 3544 8444 3596
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 9404 3544 9456 3596
rect 5540 3451 5592 3460
rect 5540 3417 5549 3451
rect 5549 3417 5583 3451
rect 5583 3417 5592 3451
rect 5540 3408 5592 3417
rect 2596 3383 2648 3392
rect 2596 3349 2605 3383
rect 2605 3349 2639 3383
rect 2639 3349 2648 3383
rect 2596 3340 2648 3349
rect 3240 3340 3292 3392
rect 8944 3451 8996 3460
rect 8944 3417 8953 3451
rect 8953 3417 8987 3451
rect 8987 3417 8996 3451
rect 8944 3408 8996 3417
rect 9220 3451 9272 3460
rect 9220 3417 9229 3451
rect 9229 3417 9263 3451
rect 9263 3417 9272 3451
rect 9220 3408 9272 3417
rect 5724 3383 5776 3392
rect 5724 3349 5749 3383
rect 5749 3349 5776 3383
rect 5724 3340 5776 3349
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 6828 3340 6880 3392
rect 8116 3340 8168 3392
rect 8392 3340 8444 3392
rect 10508 3340 10560 3392
rect 2829 3238 2881 3290
rect 2893 3238 2945 3290
rect 2957 3238 3009 3290
rect 3021 3238 3073 3290
rect 3085 3238 3137 3290
rect 5267 3238 5319 3290
rect 5331 3238 5383 3290
rect 5395 3238 5447 3290
rect 5459 3238 5511 3290
rect 5523 3238 5575 3290
rect 7705 3238 7757 3290
rect 7769 3238 7821 3290
rect 7833 3238 7885 3290
rect 7897 3238 7949 3290
rect 7961 3238 8013 3290
rect 10143 3238 10195 3290
rect 10207 3238 10259 3290
rect 10271 3238 10323 3290
rect 10335 3238 10387 3290
rect 10399 3238 10451 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 4712 3136 4764 3188
rect 5264 3136 5316 3188
rect 5724 3136 5776 3188
rect 2504 3068 2556 3120
rect 6000 3136 6052 3188
rect 6736 3136 6788 3188
rect 8944 3136 8996 3188
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2596 2932 2648 2984
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 5908 3068 5960 3120
rect 5172 3043 5224 3052
rect 4804 2932 4856 2984
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 5080 2932 5132 2984
rect 3608 2907 3660 2916
rect 3608 2873 3617 2907
rect 3617 2873 3651 2907
rect 3651 2873 3660 2907
rect 3608 2864 3660 2873
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 7012 2932 7064 2984
rect 6000 2864 6052 2916
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7748 3000 7800 3052
rect 9404 3068 9456 3120
rect 6368 2796 6420 2848
rect 7656 2932 7708 2984
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 7380 2796 7432 2848
rect 10232 2796 10284 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 848 2388 900 2440
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 9588 2252 9640 2304
rect 2829 2150 2881 2202
rect 2893 2150 2945 2202
rect 2957 2150 3009 2202
rect 3021 2150 3073 2202
rect 3085 2150 3137 2202
rect 5267 2150 5319 2202
rect 5331 2150 5383 2202
rect 5395 2150 5447 2202
rect 5459 2150 5511 2202
rect 5523 2150 5575 2202
rect 7705 2150 7757 2202
rect 7769 2150 7821 2202
rect 7833 2150 7885 2202
rect 7897 2150 7949 2202
rect 7961 2150 8013 2202
rect 10143 2150 10195 2202
rect 10207 2150 10259 2202
rect 10271 2150 10323 2202
rect 10335 2150 10387 2202
rect 10399 2150 10451 2202
<< metal2 >>
rect 3606 15328 3662 15337
rect 3606 15263 3662 15272
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1412 13394 1440 14447
rect 2169 13628 2477 13637
rect 2169 13626 2175 13628
rect 2231 13626 2255 13628
rect 2311 13626 2335 13628
rect 2391 13626 2415 13628
rect 2471 13626 2477 13628
rect 2231 13574 2233 13626
rect 2413 13574 2415 13626
rect 2169 13572 2175 13574
rect 2231 13572 2255 13574
rect 2311 13572 2335 13574
rect 2391 13572 2415 13574
rect 2471 13572 2477 13574
rect 2169 13563 2477 13572
rect 3054 13424 3110 13433
rect 1400 13388 1452 13394
rect 3054 13359 3110 13368
rect 1400 13330 1452 13336
rect 3068 13326 3096 13359
rect 3620 13326 3648 15263
rect 10414 14512 10470 14521
rect 10414 14447 10470 14456
rect 4607 13628 4915 13637
rect 4607 13626 4613 13628
rect 4669 13626 4693 13628
rect 4749 13626 4773 13628
rect 4829 13626 4853 13628
rect 4909 13626 4915 13628
rect 4669 13574 4671 13626
rect 4851 13574 4853 13626
rect 4607 13572 4613 13574
rect 4669 13572 4693 13574
rect 4749 13572 4773 13574
rect 4829 13572 4853 13574
rect 4909 13572 4915 13574
rect 4607 13563 4915 13572
rect 7045 13628 7353 13637
rect 7045 13626 7051 13628
rect 7107 13626 7131 13628
rect 7187 13626 7211 13628
rect 7267 13626 7291 13628
rect 7347 13626 7353 13628
rect 7107 13574 7109 13626
rect 7289 13574 7291 13626
rect 7045 13572 7051 13574
rect 7107 13572 7131 13574
rect 7187 13572 7211 13574
rect 7267 13572 7291 13574
rect 7347 13572 7353 13574
rect 7045 13563 7353 13572
rect 9483 13628 9791 13637
rect 9483 13626 9489 13628
rect 9545 13626 9569 13628
rect 9625 13626 9649 13628
rect 9705 13626 9729 13628
rect 9785 13626 9791 13628
rect 9545 13574 9547 13626
rect 9727 13574 9729 13626
rect 9483 13572 9489 13574
rect 9545 13572 9569 13574
rect 9625 13572 9649 13574
rect 9705 13572 9729 13574
rect 9785 13572 9791 13574
rect 9483 13563 9791 13572
rect 10428 13530 10456 14447
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 2228 13320 2280 13326
rect 3056 13320 3108 13326
rect 2228 13262 2280 13268
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 848 11144 900 11150
rect 846 11112 848 11121
rect 900 11112 902 11121
rect 846 11047 902 11056
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 860 10577 888 10610
rect 846 10568 902 10577
rect 846 10503 902 10512
rect 1412 9058 1440 13126
rect 1688 12850 1716 13262
rect 2240 12986 2268 13262
rect 2700 13258 2820 13274
rect 3056 13262 3108 13268
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 2700 13252 2832 13258
rect 2700 13246 2780 13252
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2608 12866 2636 12922
rect 2700 12889 2728 13246
rect 2780 13194 2832 13200
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 2829 13084 3137 13093
rect 2829 13082 2835 13084
rect 2891 13082 2915 13084
rect 2971 13082 2995 13084
rect 3051 13082 3075 13084
rect 3131 13082 3137 13084
rect 2891 13030 2893 13082
rect 3073 13030 3075 13082
rect 2829 13028 2835 13030
rect 2891 13028 2915 13030
rect 2971 13028 2995 13030
rect 3051 13028 3075 13030
rect 3131 13028 3137 13030
rect 2829 13019 3137 13028
rect 3252 12918 3280 13126
rect 3240 12912 3292 12918
rect 2424 12850 2636 12866
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 2412 12844 2636 12850
rect 2464 12838 2636 12844
rect 2412 12786 2464 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12170 1532 12582
rect 1688 12374 1716 12786
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 1964 12442 1992 12718
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1952 12436 2004 12442
rect 1872 12406 1952 12434
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 1688 12186 1716 12310
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1596 12158 1716 12186
rect 1596 11762 1624 12158
rect 1674 12064 1730 12073
rect 1674 11999 1730 12008
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11150 1624 11698
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1688 10674 1716 11999
rect 1872 11830 1900 12406
rect 1952 12378 2004 12384
rect 2056 12238 2084 12582
rect 2169 12540 2477 12549
rect 2169 12538 2175 12540
rect 2231 12538 2255 12540
rect 2311 12538 2335 12540
rect 2391 12538 2415 12540
rect 2471 12538 2477 12540
rect 2231 12486 2233 12538
rect 2413 12486 2415 12538
rect 2169 12484 2175 12486
rect 2231 12484 2255 12486
rect 2311 12484 2335 12486
rect 2391 12484 2415 12486
rect 2471 12484 2477 12486
rect 2169 12475 2477 12484
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1872 11150 1900 11766
rect 1964 11558 1992 12106
rect 2056 11762 2084 12174
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 2056 11082 2084 11698
rect 2424 11642 2452 12174
rect 2516 11898 2544 12718
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2424 11614 2544 11642
rect 2169 11452 2477 11461
rect 2169 11450 2175 11452
rect 2231 11450 2255 11452
rect 2311 11450 2335 11452
rect 2391 11450 2415 11452
rect 2471 11450 2477 11452
rect 2231 11398 2233 11450
rect 2413 11398 2415 11450
rect 2169 11396 2175 11398
rect 2231 11396 2255 11398
rect 2311 11396 2335 11398
rect 2391 11396 2415 11398
rect 2471 11396 2477 11398
rect 2169 11387 2477 11396
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2332 11082 2360 11222
rect 2516 11132 2544 11614
rect 2608 11354 2636 12838
rect 2686 12880 2742 12889
rect 3240 12854 3292 12860
rect 3344 12850 3372 13126
rect 2686 12815 2742 12824
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 2884 12730 2912 12786
rect 2700 12702 2912 12730
rect 2700 12374 2728 12702
rect 3344 12442 3372 12786
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 3528 12306 3556 13194
rect 5267 13084 5575 13093
rect 5267 13082 5273 13084
rect 5329 13082 5353 13084
rect 5409 13082 5433 13084
rect 5489 13082 5513 13084
rect 5569 13082 5575 13084
rect 5329 13030 5331 13082
rect 5511 13030 5513 13082
rect 5267 13028 5273 13030
rect 5329 13028 5353 13030
rect 5409 13028 5433 13030
rect 5489 13028 5513 13030
rect 5569 13028 5575 13030
rect 5267 13019 5575 13028
rect 7705 13084 8013 13093
rect 7705 13082 7711 13084
rect 7767 13082 7791 13084
rect 7847 13082 7871 13084
rect 7927 13082 7951 13084
rect 8007 13082 8013 13084
rect 7767 13030 7769 13082
rect 7949 13030 7951 13082
rect 7705 13028 7711 13030
rect 7767 13028 7791 13030
rect 7847 13028 7871 13030
rect 7927 13028 7951 13030
rect 8007 13028 8013 13030
rect 7705 13019 8013 13028
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 3240 12232 3292 12238
rect 3344 12209 3372 12242
rect 3424 12232 3476 12238
rect 3240 12174 3292 12180
rect 3330 12200 3386 12209
rect 2700 11898 2728 12174
rect 2829 11996 3137 12005
rect 2829 11994 2835 11996
rect 2891 11994 2915 11996
rect 2971 11994 2995 11996
rect 3051 11994 3075 11996
rect 3131 11994 3137 11996
rect 2891 11942 2893 11994
rect 3073 11942 3075 11994
rect 2829 11940 2835 11942
rect 2891 11940 2915 11942
rect 2971 11940 2995 11942
rect 3051 11940 3075 11942
rect 3131 11940 3137 11942
rect 2829 11931 3137 11940
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2964 11824 3016 11830
rect 2964 11766 3016 11772
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2596 11144 2648 11150
rect 2516 11104 2596 11132
rect 2596 11086 2648 11092
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 10198 1900 10406
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 1676 9988 1728 9994
rect 1676 9930 1728 9936
rect 1504 9625 1532 9930
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1412 9030 1624 9058
rect 848 8968 900 8974
rect 846 8936 848 8945
rect 1492 8968 1544 8974
rect 900 8936 902 8945
rect 1492 8910 1544 8916
rect 846 8871 902 8880
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 7993 1440 8366
rect 1398 7984 1454 7993
rect 1398 7919 1454 7928
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 848 7404 900 7410
rect 848 7346 900 7352
rect 860 7313 888 7346
rect 846 7304 902 7313
rect 846 7239 902 7248
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1412 5794 1440 7482
rect 1320 5766 1440 5794
rect 1320 5386 1348 5766
rect 1504 5710 1532 8910
rect 1596 7313 1624 9030
rect 1688 8090 1716 9930
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1780 9518 1808 9658
rect 1872 9586 1900 9862
rect 1964 9586 1992 10474
rect 2169 10364 2477 10373
rect 2169 10362 2175 10364
rect 2231 10362 2255 10364
rect 2311 10362 2335 10364
rect 2391 10362 2415 10364
rect 2471 10362 2477 10364
rect 2231 10310 2233 10362
rect 2413 10310 2415 10362
rect 2169 10308 2175 10310
rect 2231 10308 2255 10310
rect 2311 10308 2335 10310
rect 2391 10308 2415 10310
rect 2471 10308 2477 10310
rect 2169 10299 2477 10308
rect 2608 10010 2636 11086
rect 2884 11082 2912 11562
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2976 11014 3004 11766
rect 3252 11762 3280 12174
rect 3424 12174 3476 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3330 12135 3386 12144
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11150 3188 11494
rect 3252 11286 3280 11698
rect 3436 11558 3464 12174
rect 3608 12164 3660 12170
rect 3608 12106 3660 12112
rect 3620 11762 3648 12106
rect 3896 11898 3924 12174
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3988 11778 4016 12310
rect 4160 12232 4212 12238
rect 3896 11762 4016 11778
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3884 11756 4016 11762
rect 3936 11750 4016 11756
rect 4080 12192 4160 12220
rect 3884 11698 3936 11704
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3436 11354 3464 11494
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3804 11286 3832 11494
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3240 11144 3292 11150
rect 3424 11144 3476 11150
rect 3240 11086 3292 11092
rect 3344 11104 3424 11132
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2829 10908 3137 10917
rect 2829 10906 2835 10908
rect 2891 10906 2915 10908
rect 2971 10906 2995 10908
rect 3051 10906 3075 10908
rect 3131 10906 3137 10908
rect 2891 10854 2893 10906
rect 3073 10854 3075 10906
rect 2829 10852 2835 10854
rect 2891 10852 2915 10854
rect 2971 10852 2995 10854
rect 3051 10852 3075 10854
rect 3131 10852 3137 10854
rect 2829 10843 3137 10852
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2976 10062 3004 10202
rect 2872 10056 2924 10062
rect 2608 9994 2728 10010
rect 2872 9998 2924 10004
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 2608 9988 2740 9994
rect 2608 9982 2688 9988
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1964 9178 1992 9522
rect 2056 9518 2084 9930
rect 2608 9722 2636 9982
rect 2688 9930 2740 9936
rect 2884 9926 2912 9998
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2829 9820 3137 9829
rect 2829 9818 2835 9820
rect 2891 9818 2915 9820
rect 2971 9818 2995 9820
rect 3051 9818 3075 9820
rect 3131 9818 3137 9820
rect 2891 9766 2893 9818
rect 3073 9766 3075 9818
rect 2829 9764 2835 9766
rect 2891 9764 2915 9766
rect 2971 9764 2995 9766
rect 3051 9764 3075 9766
rect 3131 9764 3137 9766
rect 2829 9755 3137 9764
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2608 8974 2636 9658
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 9466 2820 9590
rect 3252 9586 3280 11086
rect 3344 10062 3372 11104
rect 3424 11086 3476 11092
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9512 3200 9518
rect 2792 9460 3148 9466
rect 2792 9454 3200 9460
rect 2792 9438 3188 9454
rect 3068 8974 3096 9438
rect 3252 9382 3280 9522
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3160 9058 3188 9318
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3160 9030 3280 9058
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1688 7410 1716 8026
rect 1780 7478 1808 8366
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1582 7304 1638 7313
rect 1582 7239 1638 7248
rect 1596 6798 1624 7239
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1688 6662 1716 7346
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1596 6458 1624 6598
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1780 6322 1808 6734
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1320 5358 1440 5386
rect 848 4616 900 4622
rect 846 4584 848 4593
rect 900 4584 902 4593
rect 846 4519 902 4528
rect 1412 4282 1440 5358
rect 1504 5234 1532 5646
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1596 5098 1624 6258
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1596 4486 1624 5034
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 4049 888 4082
rect 846 4040 902 4049
rect 846 3975 902 3984
rect 1412 3534 1440 4218
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3670 1624 3878
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 848 3460 900 3466
rect 848 3402 900 3408
rect 860 3233 888 3402
rect 846 3224 902 3233
rect 846 3159 902 3168
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 900 2408 902 2417
rect 846 2343 902 2352
rect 1504 1465 1532 2994
rect 1688 2514 1716 5170
rect 1780 3602 1808 6258
rect 1872 4826 1900 8842
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8022 2084 8774
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2056 7342 2084 7958
rect 2516 7886 2544 8910
rect 2608 8090 2636 8910
rect 2829 8732 3137 8741
rect 2829 8730 2835 8732
rect 2891 8730 2915 8732
rect 2971 8730 2995 8732
rect 3051 8730 3075 8732
rect 3131 8730 3137 8732
rect 2891 8678 2893 8730
rect 3073 8678 3075 8730
rect 2829 8676 2835 8678
rect 2891 8676 2915 8678
rect 2971 8676 2995 8678
rect 3051 8676 3075 8678
rect 3131 8676 3137 8678
rect 2829 8667 3137 8676
rect 3252 8498 3280 9030
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2608 7818 2636 8026
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2424 7206 2452 7686
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1964 6390 1992 6666
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5234 1992 6190
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1964 4214 1992 5170
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2056 3602 2084 7142
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2424 6798 2452 6870
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2240 6254 2268 6734
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2516 5778 2544 7686
rect 2608 7478 2636 7754
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2700 6934 2728 7958
rect 2829 7644 3137 7653
rect 2829 7642 2835 7644
rect 2891 7642 2915 7644
rect 2971 7642 2995 7644
rect 3051 7642 3075 7644
rect 3131 7642 3137 7644
rect 2891 7590 2893 7642
rect 3073 7590 3075 7642
rect 2829 7588 2835 7590
rect 2891 7588 2915 7590
rect 2971 7588 2995 7590
rect 3051 7588 3075 7590
rect 3131 7588 3137 7590
rect 2829 7579 3137 7588
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 7002 2820 7142
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 2976 6798 3004 6831
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2700 6202 2728 6734
rect 2829 6556 3137 6565
rect 2829 6554 2835 6556
rect 2891 6554 2915 6556
rect 2971 6554 2995 6556
rect 3051 6554 3075 6556
rect 3131 6554 3137 6556
rect 2891 6502 2893 6554
rect 3073 6502 3075 6554
rect 2829 6500 2835 6502
rect 2891 6500 2915 6502
rect 2971 6500 2995 6502
rect 3051 6500 3075 6502
rect 3131 6500 3137 6502
rect 2829 6491 3137 6500
rect 3252 6390 3280 7278
rect 3344 6458 3372 9998
rect 3528 9926 3556 11018
rect 3896 10130 3924 11698
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 10713 4016 11630
rect 4080 11014 4108 12192
rect 4160 12174 4212 12180
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11762 4200 12038
rect 4448 11830 4476 12310
rect 4436 11824 4488 11830
rect 4540 11801 4568 12582
rect 4607 12540 4915 12549
rect 4607 12538 4613 12540
rect 4669 12538 4693 12540
rect 4749 12538 4773 12540
rect 4829 12538 4853 12540
rect 4909 12538 4915 12540
rect 4669 12486 4671 12538
rect 4851 12486 4853 12538
rect 4607 12484 4613 12486
rect 4669 12484 4693 12486
rect 4749 12484 4773 12486
rect 4829 12484 4853 12486
rect 4909 12484 4915 12486
rect 4607 12475 4915 12484
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4724 11830 4752 12310
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11824 4764 11830
rect 4436 11766 4488 11772
rect 4526 11792 4582 11801
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4344 11756 4396 11762
rect 4712 11766 4764 11772
rect 4526 11727 4582 11736
rect 4344 11698 4396 11704
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4172 11354 4200 11562
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4264 11218 4292 11562
rect 4356 11286 4384 11698
rect 4816 11558 4844 12038
rect 4908 11642 4936 12242
rect 5000 11898 5028 12922
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4986 11792 5042 11801
rect 4986 11727 4988 11736
rect 5040 11727 5042 11736
rect 5092 11744 5120 12242
rect 5184 11898 5212 12718
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5552 12322 5580 12650
rect 5908 12368 5960 12374
rect 5552 12294 5764 12322
rect 6092 12368 6144 12374
rect 5908 12310 5960 12316
rect 6090 12336 6092 12345
rect 6144 12336 6146 12345
rect 5552 12238 5580 12294
rect 5540 12232 5592 12238
rect 5632 12232 5684 12238
rect 5540 12174 5592 12180
rect 5630 12200 5632 12209
rect 5684 12200 5686 12209
rect 5630 12135 5686 12144
rect 5632 12096 5684 12102
rect 5736 12073 5764 12294
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5632 12038 5684 12044
rect 5722 12064 5778 12073
rect 5267 11996 5575 12005
rect 5267 11994 5273 11996
rect 5329 11994 5353 11996
rect 5409 11994 5433 11996
rect 5489 11994 5513 11996
rect 5569 11994 5575 11996
rect 5329 11942 5331 11994
rect 5511 11942 5513 11994
rect 5267 11940 5273 11942
rect 5329 11940 5353 11942
rect 5409 11940 5433 11942
rect 5489 11940 5513 11942
rect 5569 11940 5575 11942
rect 5267 11931 5575 11940
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5644 11762 5672 12038
rect 5722 11999 5778 12008
rect 5540 11756 5592 11762
rect 5092 11716 5540 11744
rect 4988 11698 5040 11704
rect 5540 11698 5592 11704
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 4908 11614 5028 11642
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4448 11286 4476 11494
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3988 10130 4016 10202
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9110 3556 9862
rect 3988 9722 4016 10066
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4080 9654 4108 10950
rect 4172 10606 4200 11086
rect 4264 10674 4292 11154
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 9722 4200 10542
rect 4356 10470 4384 11222
rect 4540 11218 4568 11494
rect 4607 11452 4915 11461
rect 4607 11450 4613 11452
rect 4669 11450 4693 11452
rect 4749 11450 4773 11452
rect 4829 11450 4853 11452
rect 4909 11450 4915 11452
rect 4669 11398 4671 11450
rect 4851 11398 4853 11450
rect 4607 11396 4613 11398
rect 4669 11396 4693 11398
rect 4749 11396 4773 11398
rect 4829 11396 4853 11398
rect 4909 11396 4915 11398
rect 4607 11387 4915 11396
rect 5000 11354 5028 11614
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4988 11348 5040 11354
rect 5040 11308 5120 11336
rect 4988 11290 5040 11296
rect 4804 11280 4856 11286
rect 4856 11228 5028 11234
rect 4804 11222 5028 11228
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4816 11206 5028 11222
rect 4816 11150 4844 11206
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3804 9042 3832 9522
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3896 9178 3924 9454
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7410 3924 7686
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3514 6896 3570 6905
rect 3988 6866 4016 9454
rect 4080 9450 4108 9590
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4448 8922 4476 10639
rect 4264 8894 4476 8922
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3976 6860 4028 6866
rect 3514 6831 3570 6840
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3436 6322 3464 6666
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2608 6174 2728 6202
rect 2608 6118 2636 6174
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2240 5234 2268 5646
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2504 5228 2556 5234
rect 2608 5216 2636 6054
rect 2829 5468 3137 5477
rect 2829 5466 2835 5468
rect 2891 5466 2915 5468
rect 2971 5466 2995 5468
rect 3051 5466 3075 5468
rect 3131 5466 3137 5468
rect 2891 5414 2893 5466
rect 3073 5414 3075 5466
rect 2829 5412 2835 5414
rect 2891 5412 2915 5414
rect 2971 5412 2995 5414
rect 3051 5412 3075 5414
rect 3131 5412 3137 5414
rect 2829 5403 3137 5412
rect 3528 5370 3556 6831
rect 3896 6820 3976 6848
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 2884 5234 2912 5306
rect 2556 5188 2636 5216
rect 2872 5228 2924 5234
rect 2504 5170 2556 5176
rect 2872 5170 2924 5176
rect 2240 5030 2268 5170
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4146 2176 4422
rect 2516 4282 2544 5170
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 2829 4380 3137 4389
rect 2829 4378 2835 4380
rect 2891 4378 2915 4380
rect 2971 4378 2995 4380
rect 3051 4378 3075 4380
rect 3131 4378 3137 4380
rect 2891 4326 2893 4378
rect 3073 4326 3075 4378
rect 2829 4324 2835 4326
rect 2891 4324 2915 4326
rect 2971 4324 2995 4326
rect 3051 4324 3075 4326
rect 3131 4324 3137 4326
rect 2829 4315 3137 4324
rect 3436 4282 3464 4558
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3528 4214 3556 5306
rect 3804 4554 3832 5510
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3516 4208 3568 4214
rect 2318 4176 2374 4185
rect 2136 4140 2188 4146
rect 3516 4150 3568 4156
rect 3804 4146 3832 4490
rect 3896 4486 3924 6820
rect 3976 6802 4028 6808
rect 4080 6254 4108 8774
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7886 4200 8230
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7410 4200 7822
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4264 7290 4292 8894
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 7954 4384 8774
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7954 4476 8230
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4448 7546 4476 7890
rect 4540 7886 4568 11018
rect 4632 10810 4660 11086
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4908 10538 4936 11086
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4607 10364 4915 10373
rect 4607 10362 4613 10364
rect 4669 10362 4693 10364
rect 4749 10362 4773 10364
rect 4829 10362 4853 10364
rect 4909 10362 4915 10364
rect 4669 10310 4671 10362
rect 4851 10310 4853 10362
rect 4607 10308 4613 10310
rect 4669 10308 4693 10310
rect 4749 10308 4773 10310
rect 4829 10308 4853 10310
rect 4909 10308 4915 10310
rect 4607 10299 4915 10308
rect 5000 9518 5028 11206
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8362 4660 8434
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7410 4568 7822
rect 4632 7410 4660 7958
rect 4724 7954 4752 8026
rect 5000 7954 5028 8230
rect 5092 8090 5120 11308
rect 5184 10266 5212 11494
rect 5276 11218 5304 11562
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5267 10908 5575 10917
rect 5267 10906 5273 10908
rect 5329 10906 5353 10908
rect 5409 10906 5433 10908
rect 5489 10906 5513 10908
rect 5569 10906 5575 10908
rect 5329 10854 5331 10906
rect 5511 10854 5513 10906
rect 5267 10852 5273 10854
rect 5329 10852 5353 10854
rect 5409 10852 5433 10854
rect 5489 10852 5513 10854
rect 5569 10852 5575 10854
rect 5267 10843 5575 10852
rect 5736 10810 5764 11999
rect 5828 11801 5856 12242
rect 5814 11792 5870 11801
rect 5920 11762 5948 12310
rect 6090 12271 6146 12280
rect 6288 12102 6316 12718
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6090 11792 6146 11801
rect 5814 11727 5870 11736
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5920 11665 5948 11698
rect 5906 11656 5962 11665
rect 5906 11591 5962 11600
rect 6012 10810 6040 11766
rect 6090 11727 6146 11736
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5724 10804 5776 10810
rect 6000 10804 6052 10810
rect 5724 10746 5776 10752
rect 5920 10764 6000 10792
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5276 10112 5304 10746
rect 5446 10704 5502 10713
rect 5446 10639 5448 10648
rect 5500 10639 5502 10648
rect 5816 10668 5868 10674
rect 5448 10610 5500 10616
rect 5816 10610 5868 10616
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5184 10084 5304 10112
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4264 7262 4384 7290
rect 4632 7274 4660 7346
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4172 6934 4200 7142
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4264 6798 4292 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4356 6746 4384 7262
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4448 6866 4476 7210
rect 4724 7206 4752 7890
rect 5000 7546 5028 7890
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5092 7426 5120 7754
rect 5000 7410 5120 7426
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4988 7404 5120 7410
rect 5040 7398 5120 7404
rect 4988 7346 5040 7352
rect 4712 7200 4764 7206
rect 4908 7188 4936 7346
rect 5080 7200 5132 7206
rect 4908 7160 5028 7188
rect 4712 7142 4764 7148
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4620 6928 4672 6934
rect 5000 6916 5028 7160
rect 5080 7142 5132 7148
rect 4620 6870 4672 6876
rect 4816 6888 5028 6916
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4172 5370 4200 6326
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5352 4292 6734
rect 4356 6730 4476 6746
rect 4356 6724 4488 6730
rect 4356 6718 4436 6724
rect 4356 6118 4384 6718
rect 4436 6666 4488 6672
rect 4344 6112 4396 6118
rect 4632 6100 4660 6870
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 6458 4752 6734
rect 4816 6662 4844 6888
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4908 6390 4936 6734
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4632 6072 5028 6100
rect 4344 6054 4396 6060
rect 4356 5710 4384 6054
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4264 5324 4476 5352
rect 4264 5250 4292 5324
rect 4448 5284 4476 5324
rect 4528 5296 4580 5302
rect 4448 5256 4528 5284
rect 4080 5234 4292 5250
rect 4528 5238 4580 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4068 5228 4292 5234
rect 4120 5222 4292 5228
rect 4068 5170 4120 5176
rect 3988 4758 4016 5170
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 5030 4200 5102
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 4554 4016 4694
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3988 4146 4016 4490
rect 4264 4146 4292 5222
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4356 4826 4384 5170
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4448 4570 4476 4966
rect 4540 4808 4568 5238
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4540 4780 4752 4808
rect 4724 4622 4752 4780
rect 4620 4616 4672 4622
rect 4356 4564 4620 4570
rect 4356 4558 4672 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4356 4542 4660 4558
rect 4356 4146 4384 4542
rect 4816 4486 4844 4558
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4816 4282 4844 4422
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4908 4146 4936 4422
rect 2318 4111 2320 4120
rect 2136 4082 2188 4088
rect 2372 4111 2374 4120
rect 2504 4140 2556 4146
rect 2320 4082 2372 4088
rect 2504 4082 2556 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1964 3097 1992 3130
rect 2516 3126 2544 4082
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3252 3398 3280 3878
rect 3344 3534 3372 3878
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3608 3528 3660 3534
rect 3896 3505 3924 3946
rect 4448 3738 4476 4014
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4712 3664 4764 3670
rect 4710 3632 4712 3641
rect 4764 3632 4766 3641
rect 4710 3567 4766 3576
rect 4712 3528 4764 3534
rect 3608 3470 3660 3476
rect 3882 3496 3938 3505
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2504 3120 2556 3126
rect 1950 3088 2006 3097
rect 1768 3052 1820 3058
rect 2504 3062 2556 3068
rect 1950 3023 2006 3032
rect 1768 2994 1820 3000
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 1780 649 1808 2994
rect 2608 2990 2636 3334
rect 2829 3292 3137 3301
rect 2829 3290 2835 3292
rect 2891 3290 2915 3292
rect 2971 3290 2995 3292
rect 3051 3290 3075 3292
rect 3131 3290 3137 3292
rect 2891 3238 2893 3290
rect 3073 3238 3075 3290
rect 2829 3236 2835 3238
rect 2891 3236 2915 3238
rect 2971 3236 2995 3238
rect 3051 3236 3075 3238
rect 3131 3236 3137 3238
rect 2829 3227 3137 3236
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 3620 2922 3648 3470
rect 4712 3470 4764 3476
rect 3882 3431 3938 3440
rect 3896 3058 3924 3431
rect 4724 3194 4752 3470
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4804 2984 4856 2990
rect 5000 2972 5028 6072
rect 5092 5030 5120 7142
rect 5184 6882 5212 10084
rect 5460 10062 5488 10474
rect 5828 10266 5856 10610
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5267 9820 5575 9829
rect 5267 9818 5273 9820
rect 5329 9818 5353 9820
rect 5409 9818 5433 9820
rect 5489 9818 5513 9820
rect 5569 9818 5575 9820
rect 5329 9766 5331 9818
rect 5511 9766 5513 9818
rect 5267 9764 5273 9766
rect 5329 9764 5353 9766
rect 5409 9764 5433 9766
rect 5489 9764 5513 9766
rect 5569 9764 5575 9766
rect 5267 9755 5575 9764
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 8906 5396 9386
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5552 8906 5580 9046
rect 5724 8968 5776 8974
rect 5722 8936 5724 8945
rect 5776 8936 5778 8945
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5540 8900 5592 8906
rect 5722 8871 5778 8880
rect 5540 8842 5592 8848
rect 5267 8732 5575 8741
rect 5267 8730 5273 8732
rect 5329 8730 5353 8732
rect 5409 8730 5433 8732
rect 5489 8730 5513 8732
rect 5569 8730 5575 8732
rect 5329 8678 5331 8730
rect 5511 8678 5513 8730
rect 5267 8676 5273 8678
rect 5329 8676 5353 8678
rect 5409 8676 5433 8678
rect 5489 8676 5513 8678
rect 5569 8676 5575 8678
rect 5267 8667 5575 8676
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8090 5672 8230
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5267 7644 5575 7653
rect 5267 7642 5273 7644
rect 5329 7642 5353 7644
rect 5409 7642 5433 7644
rect 5489 7642 5513 7644
rect 5569 7642 5575 7644
rect 5329 7590 5331 7642
rect 5511 7590 5513 7642
rect 5267 7588 5273 7590
rect 5329 7588 5353 7590
rect 5409 7588 5433 7590
rect 5489 7588 5513 7590
rect 5569 7588 5575 7590
rect 5267 7579 5575 7588
rect 5736 7002 5764 7822
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5920 6905 5948 10764
rect 6000 10746 6052 10752
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10470 6040 10542
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10130 6040 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6000 9988 6052 9994
rect 6104 9976 6132 11727
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6196 10606 6224 11562
rect 6288 10810 6316 12038
rect 6380 11354 6408 12786
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6840 12442 6868 12582
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6932 12374 6960 12582
rect 7045 12540 7353 12549
rect 7045 12538 7051 12540
rect 7107 12538 7131 12540
rect 7187 12538 7211 12540
rect 7267 12538 7291 12540
rect 7347 12538 7353 12540
rect 7107 12486 7109 12538
rect 7289 12486 7291 12538
rect 7045 12484 7051 12486
rect 7107 12484 7131 12486
rect 7187 12484 7211 12486
rect 7267 12484 7291 12486
rect 7347 12484 7353 12486
rect 7045 12475 7353 12484
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6552 12232 6604 12238
rect 6458 12200 6514 12209
rect 6552 12174 6604 12180
rect 6458 12135 6514 12144
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6472 11257 6500 12135
rect 6564 11898 6592 12174
rect 6920 12096 6972 12102
rect 7024 12084 7052 12310
rect 7104 12232 7156 12238
rect 7102 12200 7104 12209
rect 7156 12200 7158 12209
rect 7102 12135 7158 12144
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 6972 12056 7052 12084
rect 7300 12073 7328 12106
rect 7286 12064 7342 12073
rect 6920 12038 6972 12044
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6932 11762 6960 12038
rect 7286 11999 7342 12008
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6458 11248 6514 11257
rect 6458 11183 6514 11192
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6052 9948 6132 9976
rect 6000 9930 6052 9936
rect 6012 8650 6040 9930
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 9110 6132 9454
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6104 8906 6132 9046
rect 6196 8974 6224 9522
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 8974 6316 9318
rect 6184 8968 6236 8974
rect 6182 8936 6184 8945
rect 6276 8968 6328 8974
rect 6236 8936 6238 8945
rect 6092 8900 6144 8906
rect 6276 8910 6328 8916
rect 6182 8871 6238 8880
rect 6092 8842 6144 8848
rect 6104 8786 6132 8842
rect 6104 8758 6224 8786
rect 6012 8622 6132 8650
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 8401 6040 8434
rect 5998 8392 6054 8401
rect 5998 8327 6054 8336
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7274 6040 7890
rect 6104 7449 6132 8622
rect 6090 7440 6146 7449
rect 6090 7375 6146 7384
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5906 6896 5962 6905
rect 5184 6854 5764 6882
rect 5460 6798 5488 6854
rect 5448 6792 5500 6798
rect 5262 6760 5318 6769
rect 5448 6734 5500 6740
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5262 6695 5264 6704
rect 5316 6695 5318 6704
rect 5264 6666 5316 6672
rect 5267 6556 5575 6565
rect 5267 6554 5273 6556
rect 5329 6554 5353 6556
rect 5409 6554 5433 6556
rect 5489 6554 5513 6556
rect 5569 6554 5575 6556
rect 5329 6502 5331 6554
rect 5511 6502 5513 6554
rect 5267 6500 5273 6502
rect 5329 6500 5353 6502
rect 5409 6500 5433 6502
rect 5489 6500 5513 6502
rect 5569 6500 5575 6502
rect 5267 6491 5575 6500
rect 5644 6254 5672 6734
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5736 5574 5764 6854
rect 5906 6831 5962 6840
rect 5920 6798 5948 6831
rect 5908 6792 5960 6798
rect 5814 6760 5870 6769
rect 5908 6734 5960 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5814 6695 5870 6704
rect 5828 6458 5856 6695
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6012 6186 6040 6734
rect 6104 6322 6132 7375
rect 6196 6322 6224 8758
rect 6288 8498 6316 8910
rect 6472 8650 6500 11183
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6564 10198 6592 11086
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6564 9654 6592 10134
rect 6656 9926 6684 11494
rect 6932 11336 6960 11698
rect 7024 11558 7052 11863
rect 7392 11801 7420 12718
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 11898 7512 12582
rect 7944 12434 7972 12786
rect 8588 12714 8616 13262
rect 10143 13084 10451 13093
rect 10143 13082 10149 13084
rect 10205 13082 10229 13084
rect 10285 13082 10309 13084
rect 10365 13082 10389 13084
rect 10445 13082 10451 13084
rect 10205 13030 10207 13082
rect 10387 13030 10389 13082
rect 10143 13028 10149 13030
rect 10205 13028 10229 13030
rect 10285 13028 10309 13030
rect 10365 13028 10389 13030
rect 10445 13028 10451 13030
rect 10143 13019 10451 13028
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 9483 12540 9791 12549
rect 9483 12538 9489 12540
rect 9545 12538 9569 12540
rect 9625 12538 9649 12540
rect 9705 12538 9729 12540
rect 9785 12538 9791 12540
rect 9545 12486 9547 12538
rect 9727 12486 9729 12538
rect 9483 12484 9489 12486
rect 9545 12484 9569 12486
rect 9625 12484 9649 12486
rect 9705 12484 9729 12486
rect 9785 12484 9791 12486
rect 9483 12475 9791 12484
rect 7576 12406 7972 12434
rect 7576 12238 7604 12406
rect 7944 12374 7972 12406
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7932 12368 7984 12374
rect 10244 12345 10272 12786
rect 10416 12640 10468 12646
rect 10414 12608 10416 12617
rect 10468 12608 10470 12617
rect 10414 12543 10470 12552
rect 7932 12310 7984 12316
rect 10230 12336 10286 12345
rect 7760 12238 7788 12310
rect 10230 12271 10286 12280
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7748 12232 7800 12238
rect 8116 12232 8168 12238
rect 7748 12174 7800 12180
rect 7930 12200 7986 12209
rect 7472 11892 7524 11898
rect 7576 11880 7604 12174
rect 8116 12174 8168 12180
rect 7930 12135 7932 12144
rect 7984 12135 7986 12144
rect 7932 12106 7984 12112
rect 7705 11996 8013 12005
rect 7705 11994 7711 11996
rect 7767 11994 7791 11996
rect 7847 11994 7871 11996
rect 7927 11994 7951 11996
rect 8007 11994 8013 11996
rect 7767 11942 7769 11994
rect 7949 11942 7951 11994
rect 7705 11940 7711 11942
rect 7767 11940 7791 11942
rect 7847 11940 7871 11942
rect 7927 11940 7951 11942
rect 8007 11940 8013 11942
rect 7705 11931 8013 11940
rect 7748 11892 7800 11898
rect 7576 11852 7748 11880
rect 7472 11834 7524 11840
rect 7748 11834 7800 11840
rect 7378 11792 7434 11801
rect 7196 11756 7248 11762
rect 7760 11762 7788 11834
rect 7378 11727 7434 11736
rect 7472 11756 7524 11762
rect 7196 11698 7248 11704
rect 7472 11698 7524 11704
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7208 11642 7236 11698
rect 7208 11614 7420 11642
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7045 11452 7353 11461
rect 7045 11450 7051 11452
rect 7107 11450 7131 11452
rect 7187 11450 7211 11452
rect 7267 11450 7291 11452
rect 7347 11450 7353 11452
rect 7107 11398 7109 11450
rect 7289 11398 7291 11450
rect 7045 11396 7051 11398
rect 7107 11396 7131 11398
rect 7187 11396 7211 11398
rect 7267 11396 7291 11398
rect 7347 11396 7353 11398
rect 7045 11387 7353 11396
rect 6932 11308 7236 11336
rect 6932 11218 6960 11308
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10826 7144 11018
rect 6840 10798 7144 10826
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6656 8974 6684 9862
rect 6840 9586 6868 10798
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6932 9518 6960 10610
rect 7208 10588 7236 11308
rect 7392 10742 7420 11614
rect 7484 11354 7512 11698
rect 7576 11665 7604 11698
rect 7562 11656 7618 11665
rect 7562 11591 7618 11600
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7484 10674 7512 11290
rect 7760 11082 7788 11698
rect 8128 11558 8156 12174
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8220 11812 8248 12038
rect 8300 11824 8352 11830
rect 8220 11784 8300 11812
rect 8220 11665 8248 11784
rect 8300 11766 8352 11772
rect 9324 11762 9352 12038
rect 10143 11996 10451 12005
rect 10143 11994 10149 11996
rect 10205 11994 10229 11996
rect 10285 11994 10309 11996
rect 10365 11994 10389 11996
rect 10445 11994 10451 11996
rect 10205 11942 10207 11994
rect 10387 11942 10389 11994
rect 10143 11940 10149 11942
rect 10205 11940 10229 11942
rect 10285 11940 10309 11942
rect 10365 11940 10389 11942
rect 10445 11940 10451 11942
rect 10143 11931 10451 11940
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8392 11688 8444 11694
rect 8206 11656 8262 11665
rect 8392 11630 8444 11636
rect 8206 11591 8262 11600
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7944 11286 7972 11494
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 8036 11082 8064 11290
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7705 10908 8013 10917
rect 7705 10906 7711 10908
rect 7767 10906 7791 10908
rect 7847 10906 7871 10908
rect 7927 10906 7951 10908
rect 8007 10906 8013 10908
rect 7767 10854 7769 10906
rect 7949 10854 7951 10906
rect 7705 10852 7711 10854
rect 7767 10852 7791 10854
rect 7847 10852 7871 10854
rect 7927 10852 7951 10854
rect 8007 10852 8013 10854
rect 7705 10843 8013 10852
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 8024 10600 8076 10606
rect 7208 10560 7420 10588
rect 7045 10364 7353 10373
rect 7045 10362 7051 10364
rect 7107 10362 7131 10364
rect 7187 10362 7211 10364
rect 7267 10362 7291 10364
rect 7347 10362 7353 10364
rect 7107 10310 7109 10362
rect 7289 10310 7291 10362
rect 7045 10308 7051 10310
rect 7107 10308 7131 10310
rect 7187 10308 7211 10310
rect 7267 10308 7291 10310
rect 7347 10308 7353 10310
rect 7045 10299 7353 10308
rect 6920 9512 6972 9518
rect 6748 9460 6920 9466
rect 6748 9454 6972 9460
rect 6748 9438 6960 9454
rect 6748 9110 6776 9438
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9110 6960 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6644 8968 6696 8974
rect 6564 8916 6644 8922
rect 6564 8910 6696 8916
rect 6564 8894 6684 8910
rect 6564 8838 6592 8894
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6472 8622 6592 8650
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6274 8392 6330 8401
rect 6274 8327 6330 8336
rect 6288 6798 6316 8327
rect 6472 8090 6500 8502
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6276 6792 6328 6798
rect 6274 6760 6276 6769
rect 6368 6792 6420 6798
rect 6328 6760 6330 6769
rect 6368 6734 6420 6740
rect 6274 6695 6330 6704
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5267 5468 5575 5477
rect 5267 5466 5273 5468
rect 5329 5466 5353 5468
rect 5409 5466 5433 5468
rect 5489 5466 5513 5468
rect 5569 5466 5575 5468
rect 5329 5414 5331 5466
rect 5511 5414 5513 5466
rect 5267 5412 5273 5414
rect 5329 5412 5353 5414
rect 5409 5412 5433 5414
rect 5489 5412 5513 5414
rect 5569 5412 5575 5414
rect 5267 5403 5575 5412
rect 6012 5234 6040 5782
rect 6104 5778 6132 6258
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4826 5120 4966
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5092 4214 5120 4762
rect 5920 4758 5948 5170
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5184 4078 5212 4626
rect 5267 4380 5575 4389
rect 5267 4378 5273 4380
rect 5329 4378 5353 4380
rect 5409 4378 5433 4380
rect 5489 4378 5513 4380
rect 5569 4378 5575 4380
rect 5329 4326 5331 4378
rect 5511 4326 5513 4378
rect 5267 4324 5273 4326
rect 5329 4324 5353 4326
rect 5409 4324 5433 4326
rect 5489 4324 5513 4326
rect 5569 4324 5575 4326
rect 5267 4315 5575 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3670 5120 3946
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5092 2990 5120 3606
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3058 5212 3538
rect 5460 3534 5488 3878
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5552 3466 5580 4218
rect 6196 3641 6224 6258
rect 6288 6186 6316 6695
rect 6380 6458 6408 6734
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6288 5642 6316 6122
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6564 5370 6592 8622
rect 6656 8566 6684 8774
rect 6644 8560 6696 8566
rect 6932 8514 6960 9046
rect 6644 8502 6696 8508
rect 6656 7954 6684 8502
rect 6840 8486 6960 8514
rect 6840 8430 6868 8486
rect 6828 8424 6880 8430
rect 7024 8378 7052 9114
rect 7392 9058 7420 10560
rect 8128 10588 8156 11494
rect 8404 11354 8432 11630
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9483 11452 9791 11461
rect 9483 11450 9489 11452
rect 9545 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9791 11452
rect 9545 11398 9547 11450
rect 9727 11398 9729 11450
rect 9483 11396 9489 11398
rect 9545 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9791 11398
rect 9483 11387 9791 11396
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 9126 11248 9182 11257
rect 8220 10674 8248 11222
rect 9784 11218 9812 11290
rect 9126 11183 9128 11192
rect 9180 11183 9182 11192
rect 9772 11212 9824 11218
rect 9128 11154 9180 11160
rect 9772 11154 9824 11160
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10810 9076 10950
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8076 10560 8156 10588
rect 8024 10542 8076 10548
rect 7705 9820 8013 9829
rect 7705 9818 7711 9820
rect 7767 9818 7791 9820
rect 7847 9818 7871 9820
rect 7927 9818 7951 9820
rect 8007 9818 8013 9820
rect 7767 9766 7769 9818
rect 7949 9766 7951 9818
rect 7705 9764 7711 9766
rect 7767 9764 7791 9766
rect 7847 9764 7871 9766
rect 7927 9764 7951 9766
rect 8007 9764 8013 9766
rect 7705 9755 8013 9764
rect 8128 9654 8156 10560
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7208 9030 7420 9058
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7116 8430 7144 8842
rect 7208 8838 7236 9030
rect 8036 8974 8064 9454
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7208 8514 7236 8774
rect 7300 8634 7328 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7208 8498 7328 8514
rect 7208 8492 7340 8498
rect 7208 8486 7288 8492
rect 7288 8434 7340 8440
rect 6828 8366 6880 8372
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6748 7732 6776 8298
rect 6840 7954 6868 8366
rect 6932 8350 7052 8378
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7886 6960 8350
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7392 7954 7420 8910
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 8220 8838 8248 10474
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8772 9586 8800 10134
rect 8956 10130 8984 10406
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8312 8974 8340 9386
rect 8772 9178 8800 9522
rect 8956 9518 8984 10066
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 7705 8732 8013 8741
rect 7705 8730 7711 8732
rect 7767 8730 7791 8732
rect 7847 8730 7871 8732
rect 7927 8730 7951 8732
rect 8007 8730 8013 8732
rect 7767 8678 7769 8730
rect 7949 8678 7951 8730
rect 7705 8676 7711 8678
rect 7767 8676 7791 8678
rect 7847 8676 7871 8678
rect 7927 8676 7951 8678
rect 8007 8676 8013 8678
rect 7705 8667 8013 8676
rect 8128 8650 8156 8774
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 8036 8622 8156 8650
rect 8220 8634 8248 8774
rect 8208 8628 8260 8634
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 6920 7880 6972 7886
rect 7484 7834 7512 8434
rect 8036 8430 8064 8622
rect 8208 8570 8260 8576
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 6920 7822 6972 7828
rect 7392 7806 7512 7834
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 6748 7704 6960 7732
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6182 3632 6238 3641
rect 6288 3602 6316 4082
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6182 3567 6238 3576
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6380 3534 6408 4014
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5267 3292 5575 3301
rect 5267 3290 5273 3292
rect 5329 3290 5353 3292
rect 5409 3290 5433 3292
rect 5489 3290 5513 3292
rect 5569 3290 5575 3292
rect 5329 3238 5331 3290
rect 5511 3238 5513 3290
rect 5267 3236 5273 3238
rect 5329 3236 5353 3238
rect 5409 3236 5433 3238
rect 5489 3236 5513 3238
rect 5569 3236 5575 3238
rect 5267 3227 5575 3236
rect 5736 3194 5764 3334
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5276 2990 5304 3130
rect 5920 3126 5948 3334
rect 6012 3194 6040 3334
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 4856 2944 5028 2972
rect 5080 2984 5132 2990
rect 4804 2926 4856 2932
rect 5080 2926 5132 2932
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 6012 2922 6040 3130
rect 6380 3097 6408 3470
rect 6366 3088 6422 3097
rect 6472 3074 6500 5170
rect 6564 4214 6592 5306
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4146 6684 6870
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 4146 6776 6666
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6840 5914 6868 6122
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6932 5710 6960 7704
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7392 6916 7420 7806
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7300 6888 7420 6916
rect 7300 6322 7328 6888
rect 7484 6798 7512 7686
rect 7576 6798 7604 7822
rect 7705 7644 8013 7653
rect 7705 7642 7711 7644
rect 7767 7642 7791 7644
rect 7847 7642 7871 7644
rect 7927 7642 7951 7644
rect 8007 7642 8013 7644
rect 7767 7590 7769 7642
rect 7949 7590 7951 7642
rect 7705 7588 7711 7590
rect 7767 7588 7791 7590
rect 7847 7588 7871 7590
rect 7927 7588 7951 7590
rect 8007 7588 8013 7590
rect 7705 7579 8013 7588
rect 8128 6866 8156 8298
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6458 7512 6598
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 6186 7328 6258
rect 7484 6254 7512 6394
rect 7576 6338 7604 6734
rect 7705 6556 8013 6565
rect 7705 6554 7711 6556
rect 7767 6554 7791 6556
rect 7847 6554 7871 6556
rect 7927 6554 7951 6556
rect 8007 6554 8013 6556
rect 7767 6502 7769 6554
rect 7949 6502 7951 6554
rect 7705 6500 7711 6502
rect 7767 6500 7791 6502
rect 7847 6500 7871 6502
rect 7927 6500 7951 6502
rect 8007 6500 8013 6502
rect 7705 6491 8013 6500
rect 7840 6384 7892 6390
rect 7576 6310 7696 6338
rect 7840 6326 7892 6332
rect 7668 6254 7696 6310
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7392 6118 7420 6190
rect 7852 6186 7880 6326
rect 8128 6322 8156 6802
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7944 6174 8156 6202
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 7392 5914 7420 6054
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7944 5846 7972 6174
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 4185 6960 5510
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 6918 4176 6974 4185
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6736 4140 6788 4146
rect 6918 4111 6974 4120
rect 6736 4082 6788 4088
rect 6656 3618 6684 4082
rect 6932 3720 6960 4111
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 6932 3692 7052 3720
rect 6656 3590 6868 3618
rect 7024 3602 7052 3692
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6840 3482 6868 3590
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7392 3534 7420 3878
rect 6920 3528 6972 3534
rect 6840 3476 6920 3482
rect 6840 3470 6972 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 6748 3194 6776 3470
rect 6840 3454 6960 3470
rect 6828 3392 6880 3398
rect 7484 3380 7512 5714
rect 7760 5658 7788 5782
rect 7576 5630 7788 5658
rect 7576 4146 7604 5630
rect 7705 5468 8013 5477
rect 7705 5466 7711 5468
rect 7767 5466 7791 5468
rect 7847 5466 7871 5468
rect 7927 5466 7951 5468
rect 8007 5466 8013 5468
rect 7767 5414 7769 5466
rect 7949 5414 7951 5466
rect 7705 5412 7711 5414
rect 7767 5412 7791 5414
rect 7847 5412 7871 5414
rect 7927 5412 7951 5414
rect 8007 5412 8013 5414
rect 7705 5403 8013 5412
rect 7705 4380 8013 4389
rect 7705 4378 7711 4380
rect 7767 4378 7791 4380
rect 7847 4378 7871 4380
rect 7927 4378 7951 4380
rect 8007 4378 8013 4380
rect 7767 4326 7769 4378
rect 7949 4326 7951 4378
rect 7705 4324 7711 4326
rect 7767 4324 7791 4326
rect 7847 4324 7871 4326
rect 7927 4324 7951 4326
rect 8007 4324 8013 4326
rect 7705 4315 8013 4324
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 4026 7696 4150
rect 8128 4146 8156 6174
rect 8220 5846 8248 6598
rect 8312 6118 8340 8910
rect 8944 8492 8996 8498
rect 9048 8480 9076 10746
rect 9784 10554 9812 11154
rect 9876 11082 9904 11494
rect 10244 11286 10272 11766
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 10060 10674 10088 11222
rect 10143 10908 10451 10917
rect 10143 10906 10149 10908
rect 10205 10906 10229 10908
rect 10285 10906 10309 10908
rect 10365 10906 10389 10908
rect 10445 10906 10451 10908
rect 10205 10854 10207 10906
rect 10387 10854 10389 10906
rect 10143 10852 10149 10854
rect 10205 10852 10229 10854
rect 10285 10852 10309 10854
rect 10365 10852 10389 10854
rect 10445 10852 10451 10854
rect 10143 10843 10451 10852
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10428 10713 10456 10746
rect 10414 10704 10470 10713
rect 10048 10668 10100 10674
rect 10414 10639 10470 10648
rect 10048 10610 10100 10616
rect 9784 10526 10088 10554
rect 9483 10364 9791 10373
rect 9483 10362 9489 10364
rect 9545 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9791 10364
rect 9545 10310 9547 10362
rect 9727 10310 9729 10362
rect 9483 10308 9489 10310
rect 9545 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9791 10310
rect 9483 10299 9791 10308
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9586 9720 9862
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8996 8452 9076 8480
rect 8944 8434 8996 8440
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8404 8294 8432 8327
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 9048 6934 9076 8452
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9232 6798 9260 9318
rect 9324 8974 9352 9318
rect 9416 9042 9444 9454
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 10060 9058 10088 10526
rect 10143 9820 10451 9829
rect 10143 9818 10149 9820
rect 10205 9818 10229 9820
rect 10285 9818 10309 9820
rect 10365 9818 10389 9820
rect 10445 9818 10451 9820
rect 10205 9766 10207 9818
rect 10387 9766 10389 9818
rect 10143 9764 10149 9766
rect 10205 9764 10229 9766
rect 10285 9764 10309 9766
rect 10365 9764 10389 9766
rect 10445 9764 10451 9766
rect 10143 9755 10451 9764
rect 9968 9042 10088 9058
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9968 9036 10100 9042
rect 9968 9030 10048 9036
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8498 9904 8774
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9968 7154 9996 9030
rect 10048 8978 10100 8984
rect 10520 8974 10548 11222
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 8498 10088 8842
rect 10874 8800 10930 8809
rect 10143 8732 10451 8741
rect 10874 8735 10930 8744
rect 10143 8730 10149 8732
rect 10205 8730 10229 8732
rect 10285 8730 10309 8732
rect 10365 8730 10389 8732
rect 10445 8730 10451 8732
rect 10205 8678 10207 8730
rect 10387 8678 10389 8730
rect 10143 8676 10149 8678
rect 10205 8676 10229 8678
rect 10285 8676 10309 8678
rect 10365 8676 10389 8678
rect 10445 8676 10451 8678
rect 10143 8667 10451 8676
rect 10888 8634 10916 8735
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9876 7126 9996 7154
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9508 6798 9536 6870
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9220 6792 9272 6798
rect 9496 6792 9548 6798
rect 9220 6734 9272 6740
rect 9416 6752 9496 6780
rect 8404 6458 8432 6734
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8312 5710 8340 6054
rect 8496 5710 8524 6054
rect 8680 5710 8708 6598
rect 8956 6322 8984 6734
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9232 6254 9260 6734
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8404 4078 8432 5510
rect 9324 5166 9352 5510
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 7576 3998 7696 4026
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7576 3534 7604 3998
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7668 3534 7696 3878
rect 8128 3534 8156 3878
rect 8404 3602 8432 4014
rect 9416 3602 9444 6752
rect 9876 6746 9904 7126
rect 10060 7018 10088 8434
rect 10143 7644 10451 7653
rect 10143 7642 10149 7644
rect 10205 7642 10229 7644
rect 10285 7642 10309 7644
rect 10365 7642 10389 7644
rect 10445 7642 10451 7644
rect 10205 7590 10207 7642
rect 10387 7590 10389 7642
rect 10143 7588 10149 7590
rect 10205 7588 10229 7590
rect 10285 7588 10309 7590
rect 10365 7588 10389 7590
rect 10445 7588 10451 7590
rect 10143 7579 10451 7588
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9496 6734 9548 6740
rect 9784 6718 9904 6746
rect 9968 6990 10088 7018
rect 10244 7002 10272 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10232 6996 10284 7002
rect 9784 6662 9812 6718
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9876 5710 9904 6258
rect 9968 6254 9996 6990
rect 10232 6938 10284 6944
rect 10428 6905 10456 7142
rect 10414 6896 10470 6905
rect 10414 6831 10470 6840
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6254 10088 6734
rect 10143 6556 10451 6565
rect 10143 6554 10149 6556
rect 10205 6554 10229 6556
rect 10285 6554 10309 6556
rect 10365 6554 10389 6556
rect 10445 6554 10451 6556
rect 10205 6502 10207 6554
rect 10387 6502 10389 6554
rect 10143 6500 10149 6502
rect 10205 6500 10229 6502
rect 10285 6500 10309 6502
rect 10365 6500 10389 6502
rect 10445 6500 10451 6502
rect 10143 6491 10451 6500
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9968 5710 9996 6190
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9508 5234 9536 5510
rect 10143 5468 10451 5477
rect 10143 5466 10149 5468
rect 10205 5466 10229 5468
rect 10285 5466 10309 5468
rect 10365 5466 10389 5468
rect 10445 5466 10451 5468
rect 10205 5414 10207 5466
rect 10387 5414 10389 5466
rect 10143 5412 10149 5414
rect 10205 5412 10229 5414
rect 10285 5412 10309 5414
rect 10365 5412 10389 5414
rect 10445 5412 10451 5414
rect 10143 5403 10451 5412
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 10416 5024 10468 5030
rect 10414 4992 10416 5001
rect 10468 4992 10470 5001
rect 9483 4924 9791 4933
rect 10414 4927 10470 4936
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 10143 4380 10451 4389
rect 10143 4378 10149 4380
rect 10205 4378 10229 4380
rect 10285 4378 10309 4380
rect 10365 4378 10389 4380
rect 10445 4378 10451 4380
rect 10205 4326 10207 4378
rect 10387 4326 10389 4378
rect 10143 4324 10149 4326
rect 10205 4324 10229 4326
rect 10285 4324 10309 4326
rect 10365 4324 10389 4326
rect 10445 4324 10451 4326
rect 10143 4315 10451 4324
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 9218 3496 9274 3505
rect 6828 3334 6880 3340
rect 7300 3352 7512 3380
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6642 3088 6698 3097
rect 6472 3046 6642 3074
rect 6840 3058 6868 3334
rect 7300 3058 7328 3352
rect 6366 3023 6422 3032
rect 6642 3023 6644 3032
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6380 2854 6408 3023
rect 6696 3023 6698 3032
rect 6828 3052 6880 3058
rect 6644 2994 6696 3000
rect 6828 2994 6880 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7012 2984 7064 2990
rect 7576 2972 7604 3470
rect 8944 3460 8996 3466
rect 9218 3431 9220 3440
rect 8944 3402 8996 3408
rect 9272 3431 9274 3440
rect 9220 3402 9272 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 7705 3292 8013 3301
rect 7705 3290 7711 3292
rect 7767 3290 7791 3292
rect 7847 3290 7871 3292
rect 7927 3290 7951 3292
rect 8007 3290 8013 3292
rect 7767 3238 7769 3290
rect 7949 3238 7951 3290
rect 7705 3236 7711 3238
rect 7767 3236 7791 3238
rect 7847 3236 7871 3238
rect 7927 3236 7951 3238
rect 8007 3236 8013 3238
rect 7705 3227 8013 3236
rect 8128 3126 8156 3334
rect 8116 3120 8168 3126
rect 7746 3088 7802 3097
rect 8116 3062 8168 3068
rect 8404 3058 8432 3334
rect 8956 3194 8984 3402
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9416 3126 9444 3538
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10143 3292 10451 3301
rect 10143 3290 10149 3292
rect 10205 3290 10229 3292
rect 10285 3290 10309 3292
rect 10365 3290 10389 3292
rect 10445 3290 10451 3292
rect 10205 3238 10207 3290
rect 10387 3238 10389 3290
rect 10143 3236 10149 3238
rect 10205 3236 10229 3238
rect 10285 3236 10309 3238
rect 10365 3236 10389 3238
rect 10445 3236 10451 3238
rect 10143 3227 10451 3236
rect 9404 3120 9456 3126
rect 10520 3097 10548 3334
rect 9404 3062 9456 3068
rect 10506 3088 10562 3097
rect 7746 3023 7748 3032
rect 7800 3023 7802 3032
rect 8392 3052 8444 3058
rect 7748 2994 7800 3000
rect 10506 3023 10562 3032
rect 8392 2994 8444 3000
rect 7656 2984 7708 2990
rect 7576 2944 7656 2972
rect 7064 2932 7420 2938
rect 7012 2926 7420 2932
rect 7656 2926 7708 2932
rect 7024 2910 7420 2926
rect 7392 2854 7420 2910
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 10244 2446 10272 2790
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 2829 2204 3137 2213
rect 2829 2202 2835 2204
rect 2891 2202 2915 2204
rect 2971 2202 2995 2204
rect 3051 2202 3075 2204
rect 3131 2202 3137 2204
rect 2891 2150 2893 2202
rect 3073 2150 3075 2202
rect 2829 2148 2835 2150
rect 2891 2148 2915 2150
rect 2971 2148 2995 2150
rect 3051 2148 3075 2150
rect 3131 2148 3137 2150
rect 2829 2139 3137 2148
rect 5267 2204 5575 2213
rect 5267 2202 5273 2204
rect 5329 2202 5353 2204
rect 5409 2202 5433 2204
rect 5489 2202 5513 2204
rect 5569 2202 5575 2204
rect 5329 2150 5331 2202
rect 5511 2150 5513 2202
rect 5267 2148 5273 2150
rect 5329 2148 5353 2150
rect 5409 2148 5433 2150
rect 5489 2148 5513 2150
rect 5569 2148 5575 2150
rect 5267 2139 5575 2148
rect 7705 2204 8013 2213
rect 7705 2202 7711 2204
rect 7767 2202 7791 2204
rect 7847 2202 7871 2204
rect 7927 2202 7951 2204
rect 8007 2202 8013 2204
rect 7767 2150 7769 2202
rect 7949 2150 7951 2202
rect 7705 2148 7711 2150
rect 7767 2148 7791 2150
rect 7847 2148 7871 2150
rect 7927 2148 7951 2150
rect 8007 2148 8013 2150
rect 7705 2139 8013 2148
rect 9600 1193 9628 2246
rect 10143 2204 10451 2213
rect 10143 2202 10149 2204
rect 10205 2202 10229 2204
rect 10285 2202 10309 2204
rect 10365 2202 10389 2204
rect 10445 2202 10451 2204
rect 10205 2150 10207 2202
rect 10387 2150 10389 2202
rect 10143 2148 10149 2150
rect 10205 2148 10229 2150
rect 10285 2148 10309 2150
rect 10365 2148 10389 2150
rect 10445 2148 10451 2150
rect 10143 2139 10451 2148
rect 9586 1184 9642 1193
rect 9586 1119 9642 1128
rect 1766 640 1822 649
rect 1766 575 1822 584
<< via2 >>
rect 3606 15272 3662 15328
rect 1398 14456 1454 14512
rect 2175 13626 2231 13628
rect 2255 13626 2311 13628
rect 2335 13626 2391 13628
rect 2415 13626 2471 13628
rect 2175 13574 2221 13626
rect 2221 13574 2231 13626
rect 2255 13574 2285 13626
rect 2285 13574 2297 13626
rect 2297 13574 2311 13626
rect 2335 13574 2349 13626
rect 2349 13574 2361 13626
rect 2361 13574 2391 13626
rect 2415 13574 2425 13626
rect 2425 13574 2471 13626
rect 2175 13572 2231 13574
rect 2255 13572 2311 13574
rect 2335 13572 2391 13574
rect 2415 13572 2471 13574
rect 3054 13368 3110 13424
rect 10414 14456 10470 14512
rect 4613 13626 4669 13628
rect 4693 13626 4749 13628
rect 4773 13626 4829 13628
rect 4853 13626 4909 13628
rect 4613 13574 4659 13626
rect 4659 13574 4669 13626
rect 4693 13574 4723 13626
rect 4723 13574 4735 13626
rect 4735 13574 4749 13626
rect 4773 13574 4787 13626
rect 4787 13574 4799 13626
rect 4799 13574 4829 13626
rect 4853 13574 4863 13626
rect 4863 13574 4909 13626
rect 4613 13572 4669 13574
rect 4693 13572 4749 13574
rect 4773 13572 4829 13574
rect 4853 13572 4909 13574
rect 7051 13626 7107 13628
rect 7131 13626 7187 13628
rect 7211 13626 7267 13628
rect 7291 13626 7347 13628
rect 7051 13574 7097 13626
rect 7097 13574 7107 13626
rect 7131 13574 7161 13626
rect 7161 13574 7173 13626
rect 7173 13574 7187 13626
rect 7211 13574 7225 13626
rect 7225 13574 7237 13626
rect 7237 13574 7267 13626
rect 7291 13574 7301 13626
rect 7301 13574 7347 13626
rect 7051 13572 7107 13574
rect 7131 13572 7187 13574
rect 7211 13572 7267 13574
rect 7291 13572 7347 13574
rect 9489 13626 9545 13628
rect 9569 13626 9625 13628
rect 9649 13626 9705 13628
rect 9729 13626 9785 13628
rect 9489 13574 9535 13626
rect 9535 13574 9545 13626
rect 9569 13574 9599 13626
rect 9599 13574 9611 13626
rect 9611 13574 9625 13626
rect 9649 13574 9663 13626
rect 9663 13574 9675 13626
rect 9675 13574 9705 13626
rect 9729 13574 9739 13626
rect 9739 13574 9785 13626
rect 9489 13572 9545 13574
rect 9569 13572 9625 13574
rect 9649 13572 9705 13574
rect 9729 13572 9785 13574
rect 846 11092 848 11112
rect 848 11092 900 11112
rect 900 11092 902 11112
rect 846 11056 902 11092
rect 846 10512 902 10568
rect 2835 13082 2891 13084
rect 2915 13082 2971 13084
rect 2995 13082 3051 13084
rect 3075 13082 3131 13084
rect 2835 13030 2881 13082
rect 2881 13030 2891 13082
rect 2915 13030 2945 13082
rect 2945 13030 2957 13082
rect 2957 13030 2971 13082
rect 2995 13030 3009 13082
rect 3009 13030 3021 13082
rect 3021 13030 3051 13082
rect 3075 13030 3085 13082
rect 3085 13030 3131 13082
rect 2835 13028 2891 13030
rect 2915 13028 2971 13030
rect 2995 13028 3051 13030
rect 3075 13028 3131 13030
rect 1674 12008 1730 12064
rect 2175 12538 2231 12540
rect 2255 12538 2311 12540
rect 2335 12538 2391 12540
rect 2415 12538 2471 12540
rect 2175 12486 2221 12538
rect 2221 12486 2231 12538
rect 2255 12486 2285 12538
rect 2285 12486 2297 12538
rect 2297 12486 2311 12538
rect 2335 12486 2349 12538
rect 2349 12486 2361 12538
rect 2361 12486 2391 12538
rect 2415 12486 2425 12538
rect 2425 12486 2471 12538
rect 2175 12484 2231 12486
rect 2255 12484 2311 12486
rect 2335 12484 2391 12486
rect 2415 12484 2471 12486
rect 2175 11450 2231 11452
rect 2255 11450 2311 11452
rect 2335 11450 2391 11452
rect 2415 11450 2471 11452
rect 2175 11398 2221 11450
rect 2221 11398 2231 11450
rect 2255 11398 2285 11450
rect 2285 11398 2297 11450
rect 2297 11398 2311 11450
rect 2335 11398 2349 11450
rect 2349 11398 2361 11450
rect 2361 11398 2391 11450
rect 2415 11398 2425 11450
rect 2425 11398 2471 11450
rect 2175 11396 2231 11398
rect 2255 11396 2311 11398
rect 2335 11396 2391 11398
rect 2415 11396 2471 11398
rect 2686 12824 2742 12880
rect 5273 13082 5329 13084
rect 5353 13082 5409 13084
rect 5433 13082 5489 13084
rect 5513 13082 5569 13084
rect 5273 13030 5319 13082
rect 5319 13030 5329 13082
rect 5353 13030 5383 13082
rect 5383 13030 5395 13082
rect 5395 13030 5409 13082
rect 5433 13030 5447 13082
rect 5447 13030 5459 13082
rect 5459 13030 5489 13082
rect 5513 13030 5523 13082
rect 5523 13030 5569 13082
rect 5273 13028 5329 13030
rect 5353 13028 5409 13030
rect 5433 13028 5489 13030
rect 5513 13028 5569 13030
rect 7711 13082 7767 13084
rect 7791 13082 7847 13084
rect 7871 13082 7927 13084
rect 7951 13082 8007 13084
rect 7711 13030 7757 13082
rect 7757 13030 7767 13082
rect 7791 13030 7821 13082
rect 7821 13030 7833 13082
rect 7833 13030 7847 13082
rect 7871 13030 7885 13082
rect 7885 13030 7897 13082
rect 7897 13030 7927 13082
rect 7951 13030 7961 13082
rect 7961 13030 8007 13082
rect 7711 13028 7767 13030
rect 7791 13028 7847 13030
rect 7871 13028 7927 13030
rect 7951 13028 8007 13030
rect 2835 11994 2891 11996
rect 2915 11994 2971 11996
rect 2995 11994 3051 11996
rect 3075 11994 3131 11996
rect 2835 11942 2881 11994
rect 2881 11942 2891 11994
rect 2915 11942 2945 11994
rect 2945 11942 2957 11994
rect 2957 11942 2971 11994
rect 2995 11942 3009 11994
rect 3009 11942 3021 11994
rect 3021 11942 3051 11994
rect 3075 11942 3085 11994
rect 3085 11942 3131 11994
rect 2835 11940 2891 11942
rect 2915 11940 2971 11942
rect 2995 11940 3051 11942
rect 3075 11940 3131 11942
rect 1490 9560 1546 9616
rect 846 8916 848 8936
rect 848 8916 900 8936
rect 900 8916 902 8936
rect 846 8880 902 8916
rect 1398 7928 1454 7984
rect 846 7248 902 7304
rect 846 6432 902 6488
rect 2175 10362 2231 10364
rect 2255 10362 2311 10364
rect 2335 10362 2391 10364
rect 2415 10362 2471 10364
rect 2175 10310 2221 10362
rect 2221 10310 2231 10362
rect 2255 10310 2285 10362
rect 2285 10310 2297 10362
rect 2297 10310 2311 10362
rect 2335 10310 2349 10362
rect 2349 10310 2361 10362
rect 2361 10310 2391 10362
rect 2415 10310 2425 10362
rect 2425 10310 2471 10362
rect 2175 10308 2231 10310
rect 2255 10308 2311 10310
rect 2335 10308 2391 10310
rect 2415 10308 2471 10310
rect 3330 12144 3386 12200
rect 2835 10906 2891 10908
rect 2915 10906 2971 10908
rect 2995 10906 3051 10908
rect 3075 10906 3131 10908
rect 2835 10854 2881 10906
rect 2881 10854 2891 10906
rect 2915 10854 2945 10906
rect 2945 10854 2957 10906
rect 2957 10854 2971 10906
rect 2995 10854 3009 10906
rect 3009 10854 3021 10906
rect 3021 10854 3051 10906
rect 3075 10854 3085 10906
rect 3085 10854 3131 10906
rect 2835 10852 2891 10854
rect 2915 10852 2971 10854
rect 2995 10852 3051 10854
rect 3075 10852 3131 10854
rect 2835 9818 2891 9820
rect 2915 9818 2971 9820
rect 2995 9818 3051 9820
rect 3075 9818 3131 9820
rect 2835 9766 2881 9818
rect 2881 9766 2891 9818
rect 2915 9766 2945 9818
rect 2945 9766 2957 9818
rect 2957 9766 2971 9818
rect 2995 9766 3009 9818
rect 3009 9766 3021 9818
rect 3021 9766 3051 9818
rect 3075 9766 3085 9818
rect 3085 9766 3131 9818
rect 2835 9764 2891 9766
rect 2915 9764 2971 9766
rect 2995 9764 3051 9766
rect 3075 9764 3131 9766
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 1582 7248 1638 7304
rect 1398 5480 1454 5536
rect 846 4564 848 4584
rect 848 4564 900 4584
rect 900 4564 902 4584
rect 846 4528 902 4564
rect 846 3984 902 4040
rect 846 3168 902 3224
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2835 8730 2891 8732
rect 2915 8730 2971 8732
rect 2995 8730 3051 8732
rect 3075 8730 3131 8732
rect 2835 8678 2881 8730
rect 2881 8678 2891 8730
rect 2915 8678 2945 8730
rect 2945 8678 2957 8730
rect 2957 8678 2971 8730
rect 2995 8678 3009 8730
rect 3009 8678 3021 8730
rect 3021 8678 3051 8730
rect 3075 8678 3085 8730
rect 3085 8678 3131 8730
rect 2835 8676 2891 8678
rect 2915 8676 2971 8678
rect 2995 8676 3051 8678
rect 3075 8676 3131 8678
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 2835 7642 2891 7644
rect 2915 7642 2971 7644
rect 2995 7642 3051 7644
rect 3075 7642 3131 7644
rect 2835 7590 2881 7642
rect 2881 7590 2891 7642
rect 2915 7590 2945 7642
rect 2945 7590 2957 7642
rect 2957 7590 2971 7642
rect 2995 7590 3009 7642
rect 3009 7590 3021 7642
rect 3021 7590 3051 7642
rect 3075 7590 3085 7642
rect 3085 7590 3131 7642
rect 2835 7588 2891 7590
rect 2915 7588 2971 7590
rect 2995 7588 3051 7590
rect 3075 7588 3131 7590
rect 2962 6840 3018 6896
rect 2835 6554 2891 6556
rect 2915 6554 2971 6556
rect 2995 6554 3051 6556
rect 3075 6554 3131 6556
rect 2835 6502 2881 6554
rect 2881 6502 2891 6554
rect 2915 6502 2945 6554
rect 2945 6502 2957 6554
rect 2957 6502 2971 6554
rect 2995 6502 3009 6554
rect 3009 6502 3021 6554
rect 3021 6502 3051 6554
rect 3075 6502 3085 6554
rect 3085 6502 3131 6554
rect 2835 6500 2891 6502
rect 2915 6500 2971 6502
rect 2995 6500 3051 6502
rect 3075 6500 3131 6502
rect 4613 12538 4669 12540
rect 4693 12538 4749 12540
rect 4773 12538 4829 12540
rect 4853 12538 4909 12540
rect 4613 12486 4659 12538
rect 4659 12486 4669 12538
rect 4693 12486 4723 12538
rect 4723 12486 4735 12538
rect 4735 12486 4749 12538
rect 4773 12486 4787 12538
rect 4787 12486 4799 12538
rect 4799 12486 4829 12538
rect 4853 12486 4863 12538
rect 4863 12486 4909 12538
rect 4613 12484 4669 12486
rect 4693 12484 4749 12486
rect 4773 12484 4829 12486
rect 4853 12484 4909 12486
rect 4526 11736 4582 11792
rect 4986 11756 5042 11792
rect 4986 11736 4988 11756
rect 4988 11736 5040 11756
rect 5040 11736 5042 11756
rect 6090 12316 6092 12336
rect 6092 12316 6144 12336
rect 6144 12316 6146 12336
rect 5630 12180 5632 12200
rect 5632 12180 5684 12200
rect 5684 12180 5686 12200
rect 5630 12144 5686 12180
rect 5273 11994 5329 11996
rect 5353 11994 5409 11996
rect 5433 11994 5489 11996
rect 5513 11994 5569 11996
rect 5273 11942 5319 11994
rect 5319 11942 5329 11994
rect 5353 11942 5383 11994
rect 5383 11942 5395 11994
rect 5395 11942 5409 11994
rect 5433 11942 5447 11994
rect 5447 11942 5459 11994
rect 5459 11942 5489 11994
rect 5513 11942 5523 11994
rect 5523 11942 5569 11994
rect 5273 11940 5329 11942
rect 5353 11940 5409 11942
rect 5433 11940 5489 11942
rect 5513 11940 5569 11942
rect 5722 12008 5778 12064
rect 3974 10648 4030 10704
rect 4613 11450 4669 11452
rect 4693 11450 4749 11452
rect 4773 11450 4829 11452
rect 4853 11450 4909 11452
rect 4613 11398 4659 11450
rect 4659 11398 4669 11450
rect 4693 11398 4723 11450
rect 4723 11398 4735 11450
rect 4735 11398 4749 11450
rect 4773 11398 4787 11450
rect 4787 11398 4799 11450
rect 4799 11398 4829 11450
rect 4853 11398 4863 11450
rect 4863 11398 4909 11450
rect 4613 11396 4669 11398
rect 4693 11396 4749 11398
rect 4773 11396 4829 11398
rect 4853 11396 4909 11398
rect 4434 10648 4490 10704
rect 3514 6840 3570 6896
rect 2835 5466 2891 5468
rect 2915 5466 2971 5468
rect 2995 5466 3051 5468
rect 3075 5466 3131 5468
rect 2835 5414 2881 5466
rect 2881 5414 2891 5466
rect 2915 5414 2945 5466
rect 2945 5414 2957 5466
rect 2957 5414 2971 5466
rect 2995 5414 3009 5466
rect 3009 5414 3021 5466
rect 3021 5414 3051 5466
rect 3075 5414 3085 5466
rect 3085 5414 3131 5466
rect 2835 5412 2891 5414
rect 2915 5412 2971 5414
rect 2995 5412 3051 5414
rect 3075 5412 3131 5414
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2835 4378 2891 4380
rect 2915 4378 2971 4380
rect 2995 4378 3051 4380
rect 3075 4378 3131 4380
rect 2835 4326 2881 4378
rect 2881 4326 2891 4378
rect 2915 4326 2945 4378
rect 2945 4326 2957 4378
rect 2957 4326 2971 4378
rect 2995 4326 3009 4378
rect 3009 4326 3021 4378
rect 3021 4326 3051 4378
rect 3075 4326 3085 4378
rect 3085 4326 3131 4378
rect 2835 4324 2891 4326
rect 2915 4324 2971 4326
rect 2995 4324 3051 4326
rect 3075 4324 3131 4326
rect 2318 4140 2374 4176
rect 4613 10362 4669 10364
rect 4693 10362 4749 10364
rect 4773 10362 4829 10364
rect 4853 10362 4909 10364
rect 4613 10310 4659 10362
rect 4659 10310 4669 10362
rect 4693 10310 4723 10362
rect 4723 10310 4735 10362
rect 4735 10310 4749 10362
rect 4773 10310 4787 10362
rect 4787 10310 4799 10362
rect 4799 10310 4829 10362
rect 4853 10310 4863 10362
rect 4863 10310 4909 10362
rect 4613 10308 4669 10310
rect 4693 10308 4749 10310
rect 4773 10308 4829 10310
rect 4853 10308 4909 10310
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 5273 10906 5329 10908
rect 5353 10906 5409 10908
rect 5433 10906 5489 10908
rect 5513 10906 5569 10908
rect 5273 10854 5319 10906
rect 5319 10854 5329 10906
rect 5353 10854 5383 10906
rect 5383 10854 5395 10906
rect 5395 10854 5409 10906
rect 5433 10854 5447 10906
rect 5447 10854 5459 10906
rect 5459 10854 5489 10906
rect 5513 10854 5523 10906
rect 5523 10854 5569 10906
rect 5273 10852 5329 10854
rect 5353 10852 5409 10854
rect 5433 10852 5489 10854
rect 5513 10852 5569 10854
rect 5814 11736 5870 11792
rect 6090 12280 6146 12316
rect 5906 11600 5962 11656
rect 6090 11736 6146 11792
rect 5446 10668 5502 10704
rect 5446 10648 5448 10668
rect 5448 10648 5500 10668
rect 5500 10648 5502 10668
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 2318 4120 2320 4140
rect 2320 4120 2372 4140
rect 2372 4120 2374 4140
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4710 3612 4712 3632
rect 4712 3612 4764 3632
rect 4764 3612 4766 3632
rect 4710 3576 4766 3612
rect 1950 3032 2006 3088
rect 1490 1400 1546 1456
rect 2835 3290 2891 3292
rect 2915 3290 2971 3292
rect 2995 3290 3051 3292
rect 3075 3290 3131 3292
rect 2835 3238 2881 3290
rect 2881 3238 2891 3290
rect 2915 3238 2945 3290
rect 2945 3238 2957 3290
rect 2957 3238 2971 3290
rect 2995 3238 3009 3290
rect 3009 3238 3021 3290
rect 3021 3238 3051 3290
rect 3075 3238 3085 3290
rect 3085 3238 3131 3290
rect 2835 3236 2891 3238
rect 2915 3236 2971 3238
rect 2995 3236 3051 3238
rect 3075 3236 3131 3238
rect 3882 3440 3938 3496
rect 5273 9818 5329 9820
rect 5353 9818 5409 9820
rect 5433 9818 5489 9820
rect 5513 9818 5569 9820
rect 5273 9766 5319 9818
rect 5319 9766 5329 9818
rect 5353 9766 5383 9818
rect 5383 9766 5395 9818
rect 5395 9766 5409 9818
rect 5433 9766 5447 9818
rect 5447 9766 5459 9818
rect 5459 9766 5489 9818
rect 5513 9766 5523 9818
rect 5523 9766 5569 9818
rect 5273 9764 5329 9766
rect 5353 9764 5409 9766
rect 5433 9764 5489 9766
rect 5513 9764 5569 9766
rect 5722 8916 5724 8936
rect 5724 8916 5776 8936
rect 5776 8916 5778 8936
rect 5722 8880 5778 8916
rect 5273 8730 5329 8732
rect 5353 8730 5409 8732
rect 5433 8730 5489 8732
rect 5513 8730 5569 8732
rect 5273 8678 5319 8730
rect 5319 8678 5329 8730
rect 5353 8678 5383 8730
rect 5383 8678 5395 8730
rect 5395 8678 5409 8730
rect 5433 8678 5447 8730
rect 5447 8678 5459 8730
rect 5459 8678 5489 8730
rect 5513 8678 5523 8730
rect 5523 8678 5569 8730
rect 5273 8676 5329 8678
rect 5353 8676 5409 8678
rect 5433 8676 5489 8678
rect 5513 8676 5569 8678
rect 5273 7642 5329 7644
rect 5353 7642 5409 7644
rect 5433 7642 5489 7644
rect 5513 7642 5569 7644
rect 5273 7590 5319 7642
rect 5319 7590 5329 7642
rect 5353 7590 5383 7642
rect 5383 7590 5395 7642
rect 5395 7590 5409 7642
rect 5433 7590 5447 7642
rect 5447 7590 5459 7642
rect 5459 7590 5489 7642
rect 5513 7590 5523 7642
rect 5523 7590 5569 7642
rect 5273 7588 5329 7590
rect 5353 7588 5409 7590
rect 5433 7588 5489 7590
rect 5513 7588 5569 7590
rect 7051 12538 7107 12540
rect 7131 12538 7187 12540
rect 7211 12538 7267 12540
rect 7291 12538 7347 12540
rect 7051 12486 7097 12538
rect 7097 12486 7107 12538
rect 7131 12486 7161 12538
rect 7161 12486 7173 12538
rect 7173 12486 7187 12538
rect 7211 12486 7225 12538
rect 7225 12486 7237 12538
rect 7237 12486 7267 12538
rect 7291 12486 7301 12538
rect 7301 12486 7347 12538
rect 7051 12484 7107 12486
rect 7131 12484 7187 12486
rect 7211 12484 7267 12486
rect 7291 12484 7347 12486
rect 6458 12144 6514 12200
rect 7102 12180 7104 12200
rect 7104 12180 7156 12200
rect 7156 12180 7158 12200
rect 7102 12144 7158 12180
rect 7286 12008 7342 12064
rect 7010 11872 7066 11928
rect 6458 11192 6514 11248
rect 6182 8916 6184 8936
rect 6184 8916 6236 8936
rect 6236 8916 6238 8936
rect 6182 8880 6238 8916
rect 5998 8336 6054 8392
rect 6090 7384 6146 7440
rect 5262 6724 5318 6760
rect 5262 6704 5264 6724
rect 5264 6704 5316 6724
rect 5316 6704 5318 6724
rect 5273 6554 5329 6556
rect 5353 6554 5409 6556
rect 5433 6554 5489 6556
rect 5513 6554 5569 6556
rect 5273 6502 5319 6554
rect 5319 6502 5329 6554
rect 5353 6502 5383 6554
rect 5383 6502 5395 6554
rect 5395 6502 5409 6554
rect 5433 6502 5447 6554
rect 5447 6502 5459 6554
rect 5459 6502 5489 6554
rect 5513 6502 5523 6554
rect 5523 6502 5569 6554
rect 5273 6500 5329 6502
rect 5353 6500 5409 6502
rect 5433 6500 5489 6502
rect 5513 6500 5569 6502
rect 5906 6840 5962 6896
rect 5814 6704 5870 6760
rect 10149 13082 10205 13084
rect 10229 13082 10285 13084
rect 10309 13082 10365 13084
rect 10389 13082 10445 13084
rect 10149 13030 10195 13082
rect 10195 13030 10205 13082
rect 10229 13030 10259 13082
rect 10259 13030 10271 13082
rect 10271 13030 10285 13082
rect 10309 13030 10323 13082
rect 10323 13030 10335 13082
rect 10335 13030 10365 13082
rect 10389 13030 10399 13082
rect 10399 13030 10445 13082
rect 10149 13028 10205 13030
rect 10229 13028 10285 13030
rect 10309 13028 10365 13030
rect 10389 13028 10445 13030
rect 9489 12538 9545 12540
rect 9569 12538 9625 12540
rect 9649 12538 9705 12540
rect 9729 12538 9785 12540
rect 9489 12486 9535 12538
rect 9535 12486 9545 12538
rect 9569 12486 9599 12538
rect 9599 12486 9611 12538
rect 9611 12486 9625 12538
rect 9649 12486 9663 12538
rect 9663 12486 9675 12538
rect 9675 12486 9705 12538
rect 9729 12486 9739 12538
rect 9739 12486 9785 12538
rect 9489 12484 9545 12486
rect 9569 12484 9625 12486
rect 9649 12484 9705 12486
rect 9729 12484 9785 12486
rect 10414 12588 10416 12608
rect 10416 12588 10468 12608
rect 10468 12588 10470 12608
rect 10414 12552 10470 12588
rect 10230 12280 10286 12336
rect 7930 12164 7986 12200
rect 7930 12144 7932 12164
rect 7932 12144 7984 12164
rect 7984 12144 7986 12164
rect 7711 11994 7767 11996
rect 7791 11994 7847 11996
rect 7871 11994 7927 11996
rect 7951 11994 8007 11996
rect 7711 11942 7757 11994
rect 7757 11942 7767 11994
rect 7791 11942 7821 11994
rect 7821 11942 7833 11994
rect 7833 11942 7847 11994
rect 7871 11942 7885 11994
rect 7885 11942 7897 11994
rect 7897 11942 7927 11994
rect 7951 11942 7961 11994
rect 7961 11942 8007 11994
rect 7711 11940 7767 11942
rect 7791 11940 7847 11942
rect 7871 11940 7927 11942
rect 7951 11940 8007 11942
rect 7378 11736 7434 11792
rect 7051 11450 7107 11452
rect 7131 11450 7187 11452
rect 7211 11450 7267 11452
rect 7291 11450 7347 11452
rect 7051 11398 7097 11450
rect 7097 11398 7107 11450
rect 7131 11398 7161 11450
rect 7161 11398 7173 11450
rect 7173 11398 7187 11450
rect 7211 11398 7225 11450
rect 7225 11398 7237 11450
rect 7237 11398 7267 11450
rect 7291 11398 7301 11450
rect 7301 11398 7347 11450
rect 7051 11396 7107 11398
rect 7131 11396 7187 11398
rect 7211 11396 7267 11398
rect 7291 11396 7347 11398
rect 7562 11600 7618 11656
rect 10149 11994 10205 11996
rect 10229 11994 10285 11996
rect 10309 11994 10365 11996
rect 10389 11994 10445 11996
rect 10149 11942 10195 11994
rect 10195 11942 10205 11994
rect 10229 11942 10259 11994
rect 10259 11942 10271 11994
rect 10271 11942 10285 11994
rect 10309 11942 10323 11994
rect 10323 11942 10335 11994
rect 10335 11942 10365 11994
rect 10389 11942 10399 11994
rect 10399 11942 10445 11994
rect 10149 11940 10205 11942
rect 10229 11940 10285 11942
rect 10309 11940 10365 11942
rect 10389 11940 10445 11942
rect 8206 11600 8262 11656
rect 7711 10906 7767 10908
rect 7791 10906 7847 10908
rect 7871 10906 7927 10908
rect 7951 10906 8007 10908
rect 7711 10854 7757 10906
rect 7757 10854 7767 10906
rect 7791 10854 7821 10906
rect 7821 10854 7833 10906
rect 7833 10854 7847 10906
rect 7871 10854 7885 10906
rect 7885 10854 7897 10906
rect 7897 10854 7927 10906
rect 7951 10854 7961 10906
rect 7961 10854 8007 10906
rect 7711 10852 7767 10854
rect 7791 10852 7847 10854
rect 7871 10852 7927 10854
rect 7951 10852 8007 10854
rect 7051 10362 7107 10364
rect 7131 10362 7187 10364
rect 7211 10362 7267 10364
rect 7291 10362 7347 10364
rect 7051 10310 7097 10362
rect 7097 10310 7107 10362
rect 7131 10310 7161 10362
rect 7161 10310 7173 10362
rect 7173 10310 7187 10362
rect 7211 10310 7225 10362
rect 7225 10310 7237 10362
rect 7237 10310 7267 10362
rect 7291 10310 7301 10362
rect 7301 10310 7347 10362
rect 7051 10308 7107 10310
rect 7131 10308 7187 10310
rect 7211 10308 7267 10310
rect 7291 10308 7347 10310
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 6274 8336 6330 8392
rect 6274 6740 6276 6760
rect 6276 6740 6328 6760
rect 6328 6740 6330 6760
rect 6274 6704 6330 6740
rect 5273 5466 5329 5468
rect 5353 5466 5409 5468
rect 5433 5466 5489 5468
rect 5513 5466 5569 5468
rect 5273 5414 5319 5466
rect 5319 5414 5329 5466
rect 5353 5414 5383 5466
rect 5383 5414 5395 5466
rect 5395 5414 5409 5466
rect 5433 5414 5447 5466
rect 5447 5414 5459 5466
rect 5459 5414 5489 5466
rect 5513 5414 5523 5466
rect 5523 5414 5569 5466
rect 5273 5412 5329 5414
rect 5353 5412 5409 5414
rect 5433 5412 5489 5414
rect 5513 5412 5569 5414
rect 5273 4378 5329 4380
rect 5353 4378 5409 4380
rect 5433 4378 5489 4380
rect 5513 4378 5569 4380
rect 5273 4326 5319 4378
rect 5319 4326 5329 4378
rect 5353 4326 5383 4378
rect 5383 4326 5395 4378
rect 5395 4326 5409 4378
rect 5433 4326 5447 4378
rect 5447 4326 5459 4378
rect 5459 4326 5489 4378
rect 5513 4326 5523 4378
rect 5523 4326 5569 4378
rect 5273 4324 5329 4326
rect 5353 4324 5409 4326
rect 5433 4324 5489 4326
rect 5513 4324 5569 4326
rect 9489 11450 9545 11452
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9489 11398 9535 11450
rect 9535 11398 9545 11450
rect 9569 11398 9599 11450
rect 9599 11398 9611 11450
rect 9611 11398 9625 11450
rect 9649 11398 9663 11450
rect 9663 11398 9675 11450
rect 9675 11398 9705 11450
rect 9729 11398 9739 11450
rect 9739 11398 9785 11450
rect 9489 11396 9545 11398
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 9126 11212 9182 11248
rect 9126 11192 9128 11212
rect 9128 11192 9180 11212
rect 9180 11192 9182 11212
rect 7711 9818 7767 9820
rect 7791 9818 7847 9820
rect 7871 9818 7927 9820
rect 7951 9818 8007 9820
rect 7711 9766 7757 9818
rect 7757 9766 7767 9818
rect 7791 9766 7821 9818
rect 7821 9766 7833 9818
rect 7833 9766 7847 9818
rect 7871 9766 7885 9818
rect 7885 9766 7897 9818
rect 7897 9766 7927 9818
rect 7951 9766 7961 9818
rect 7961 9766 8007 9818
rect 7711 9764 7767 9766
rect 7791 9764 7847 9766
rect 7871 9764 7927 9766
rect 7951 9764 8007 9766
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7711 8730 7767 8732
rect 7791 8730 7847 8732
rect 7871 8730 7927 8732
rect 7951 8730 8007 8732
rect 7711 8678 7757 8730
rect 7757 8678 7767 8730
rect 7791 8678 7821 8730
rect 7821 8678 7833 8730
rect 7833 8678 7847 8730
rect 7871 8678 7885 8730
rect 7885 8678 7897 8730
rect 7897 8678 7927 8730
rect 7951 8678 7961 8730
rect 7961 8678 8007 8730
rect 7711 8676 7767 8678
rect 7791 8676 7847 8678
rect 7871 8676 7927 8678
rect 7951 8676 8007 8678
rect 6182 3576 6238 3632
rect 5273 3290 5329 3292
rect 5353 3290 5409 3292
rect 5433 3290 5489 3292
rect 5513 3290 5569 3292
rect 5273 3238 5319 3290
rect 5319 3238 5329 3290
rect 5353 3238 5383 3290
rect 5383 3238 5395 3290
rect 5395 3238 5409 3290
rect 5433 3238 5447 3290
rect 5447 3238 5459 3290
rect 5459 3238 5489 3290
rect 5513 3238 5523 3290
rect 5523 3238 5569 3290
rect 5273 3236 5329 3238
rect 5353 3236 5409 3238
rect 5433 3236 5489 3238
rect 5513 3236 5569 3238
rect 6366 3032 6422 3088
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7711 7642 7767 7644
rect 7791 7642 7847 7644
rect 7871 7642 7927 7644
rect 7951 7642 8007 7644
rect 7711 7590 7757 7642
rect 7757 7590 7767 7642
rect 7791 7590 7821 7642
rect 7821 7590 7833 7642
rect 7833 7590 7847 7642
rect 7871 7590 7885 7642
rect 7885 7590 7897 7642
rect 7897 7590 7927 7642
rect 7951 7590 7961 7642
rect 7961 7590 8007 7642
rect 7711 7588 7767 7590
rect 7791 7588 7847 7590
rect 7871 7588 7927 7590
rect 7951 7588 8007 7590
rect 7711 6554 7767 6556
rect 7791 6554 7847 6556
rect 7871 6554 7927 6556
rect 7951 6554 8007 6556
rect 7711 6502 7757 6554
rect 7757 6502 7767 6554
rect 7791 6502 7821 6554
rect 7821 6502 7833 6554
rect 7833 6502 7847 6554
rect 7871 6502 7885 6554
rect 7885 6502 7897 6554
rect 7897 6502 7927 6554
rect 7951 6502 7961 6554
rect 7961 6502 8007 6554
rect 7711 6500 7767 6502
rect 7791 6500 7847 6502
rect 7871 6500 7927 6502
rect 7951 6500 8007 6502
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 6918 4120 6974 4176
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7711 5466 7767 5468
rect 7791 5466 7847 5468
rect 7871 5466 7927 5468
rect 7951 5466 8007 5468
rect 7711 5414 7757 5466
rect 7757 5414 7767 5466
rect 7791 5414 7821 5466
rect 7821 5414 7833 5466
rect 7833 5414 7847 5466
rect 7871 5414 7885 5466
rect 7885 5414 7897 5466
rect 7897 5414 7927 5466
rect 7951 5414 7961 5466
rect 7961 5414 8007 5466
rect 7711 5412 7767 5414
rect 7791 5412 7847 5414
rect 7871 5412 7927 5414
rect 7951 5412 8007 5414
rect 7711 4378 7767 4380
rect 7791 4378 7847 4380
rect 7871 4378 7927 4380
rect 7951 4378 8007 4380
rect 7711 4326 7757 4378
rect 7757 4326 7767 4378
rect 7791 4326 7821 4378
rect 7821 4326 7833 4378
rect 7833 4326 7847 4378
rect 7871 4326 7885 4378
rect 7885 4326 7897 4378
rect 7897 4326 7927 4378
rect 7951 4326 7961 4378
rect 7961 4326 8007 4378
rect 7711 4324 7767 4326
rect 7791 4324 7847 4326
rect 7871 4324 7927 4326
rect 7951 4324 8007 4326
rect 10149 10906 10205 10908
rect 10229 10906 10285 10908
rect 10309 10906 10365 10908
rect 10389 10906 10445 10908
rect 10149 10854 10195 10906
rect 10195 10854 10205 10906
rect 10229 10854 10259 10906
rect 10259 10854 10271 10906
rect 10271 10854 10285 10906
rect 10309 10854 10323 10906
rect 10323 10854 10335 10906
rect 10335 10854 10365 10906
rect 10389 10854 10399 10906
rect 10399 10854 10445 10906
rect 10149 10852 10205 10854
rect 10229 10852 10285 10854
rect 10309 10852 10365 10854
rect 10389 10852 10445 10854
rect 10414 10648 10470 10704
rect 9489 10362 9545 10364
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9489 10310 9535 10362
rect 9535 10310 9545 10362
rect 9569 10310 9599 10362
rect 9599 10310 9611 10362
rect 9611 10310 9625 10362
rect 9649 10310 9663 10362
rect 9663 10310 9675 10362
rect 9675 10310 9705 10362
rect 9729 10310 9739 10362
rect 9739 10310 9785 10362
rect 9489 10308 9545 10310
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 8390 8336 8446 8392
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10149 9818 10205 9820
rect 10229 9818 10285 9820
rect 10309 9818 10365 9820
rect 10389 9818 10445 9820
rect 10149 9766 10195 9818
rect 10195 9766 10205 9818
rect 10229 9766 10259 9818
rect 10259 9766 10271 9818
rect 10271 9766 10285 9818
rect 10309 9766 10323 9818
rect 10323 9766 10335 9818
rect 10335 9766 10365 9818
rect 10389 9766 10399 9818
rect 10399 9766 10445 9818
rect 10149 9764 10205 9766
rect 10229 9764 10285 9766
rect 10309 9764 10365 9766
rect 10389 9764 10445 9766
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10874 8744 10930 8800
rect 10149 8730 10205 8732
rect 10229 8730 10285 8732
rect 10309 8730 10365 8732
rect 10389 8730 10445 8732
rect 10149 8678 10195 8730
rect 10195 8678 10205 8730
rect 10229 8678 10259 8730
rect 10259 8678 10271 8730
rect 10271 8678 10285 8730
rect 10309 8678 10323 8730
rect 10323 8678 10335 8730
rect 10335 8678 10365 8730
rect 10389 8678 10399 8730
rect 10399 8678 10445 8730
rect 10149 8676 10205 8678
rect 10229 8676 10285 8678
rect 10309 8676 10365 8678
rect 10389 8676 10445 8678
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10149 7642 10205 7644
rect 10229 7642 10285 7644
rect 10309 7642 10365 7644
rect 10389 7642 10445 7644
rect 10149 7590 10195 7642
rect 10195 7590 10205 7642
rect 10229 7590 10259 7642
rect 10259 7590 10271 7642
rect 10271 7590 10285 7642
rect 10309 7590 10323 7642
rect 10323 7590 10335 7642
rect 10335 7590 10365 7642
rect 10389 7590 10399 7642
rect 10399 7590 10445 7642
rect 10149 7588 10205 7590
rect 10229 7588 10285 7590
rect 10309 7588 10365 7590
rect 10389 7588 10445 7590
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 10414 6840 10470 6896
rect 10149 6554 10205 6556
rect 10229 6554 10285 6556
rect 10309 6554 10365 6556
rect 10389 6554 10445 6556
rect 10149 6502 10195 6554
rect 10195 6502 10205 6554
rect 10229 6502 10259 6554
rect 10259 6502 10271 6554
rect 10271 6502 10285 6554
rect 10309 6502 10323 6554
rect 10323 6502 10335 6554
rect 10335 6502 10365 6554
rect 10389 6502 10399 6554
rect 10399 6502 10445 6554
rect 10149 6500 10205 6502
rect 10229 6500 10285 6502
rect 10309 6500 10365 6502
rect 10389 6500 10445 6502
rect 10149 5466 10205 5468
rect 10229 5466 10285 5468
rect 10309 5466 10365 5468
rect 10389 5466 10445 5468
rect 10149 5414 10195 5466
rect 10195 5414 10205 5466
rect 10229 5414 10259 5466
rect 10259 5414 10271 5466
rect 10271 5414 10285 5466
rect 10309 5414 10323 5466
rect 10323 5414 10335 5466
rect 10335 5414 10365 5466
rect 10389 5414 10399 5466
rect 10399 5414 10445 5466
rect 10149 5412 10205 5414
rect 10229 5412 10285 5414
rect 10309 5412 10365 5414
rect 10389 5412 10445 5414
rect 10414 4972 10416 4992
rect 10416 4972 10468 4992
rect 10468 4972 10470 4992
rect 10414 4936 10470 4972
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 10149 4378 10205 4380
rect 10229 4378 10285 4380
rect 10309 4378 10365 4380
rect 10389 4378 10445 4380
rect 10149 4326 10195 4378
rect 10195 4326 10205 4378
rect 10229 4326 10259 4378
rect 10259 4326 10271 4378
rect 10271 4326 10285 4378
rect 10309 4326 10323 4378
rect 10323 4326 10335 4378
rect 10335 4326 10365 4378
rect 10389 4326 10399 4378
rect 10399 4326 10445 4378
rect 10149 4324 10205 4326
rect 10229 4324 10285 4326
rect 10309 4324 10365 4326
rect 10389 4324 10445 4326
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 6642 3052 6698 3088
rect 6642 3032 6644 3052
rect 6644 3032 6696 3052
rect 6696 3032 6698 3052
rect 9218 3460 9274 3496
rect 9218 3440 9220 3460
rect 9220 3440 9272 3460
rect 9272 3440 9274 3460
rect 7711 3290 7767 3292
rect 7791 3290 7847 3292
rect 7871 3290 7927 3292
rect 7951 3290 8007 3292
rect 7711 3238 7757 3290
rect 7757 3238 7767 3290
rect 7791 3238 7821 3290
rect 7821 3238 7833 3290
rect 7833 3238 7847 3290
rect 7871 3238 7885 3290
rect 7885 3238 7897 3290
rect 7897 3238 7927 3290
rect 7951 3238 7961 3290
rect 7961 3238 8007 3290
rect 7711 3236 7767 3238
rect 7791 3236 7847 3238
rect 7871 3236 7927 3238
rect 7951 3236 8007 3238
rect 7746 3052 7802 3088
rect 10149 3290 10205 3292
rect 10229 3290 10285 3292
rect 10309 3290 10365 3292
rect 10389 3290 10445 3292
rect 10149 3238 10195 3290
rect 10195 3238 10205 3290
rect 10229 3238 10259 3290
rect 10259 3238 10271 3290
rect 10271 3238 10285 3290
rect 10309 3238 10323 3290
rect 10323 3238 10335 3290
rect 10335 3238 10365 3290
rect 10389 3238 10399 3290
rect 10399 3238 10445 3290
rect 10149 3236 10205 3238
rect 10229 3236 10285 3238
rect 10309 3236 10365 3238
rect 10389 3236 10445 3238
rect 7746 3032 7748 3052
rect 7748 3032 7800 3052
rect 7800 3032 7802 3052
rect 10506 3032 10562 3088
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 2835 2202 2891 2204
rect 2915 2202 2971 2204
rect 2995 2202 3051 2204
rect 3075 2202 3131 2204
rect 2835 2150 2881 2202
rect 2881 2150 2891 2202
rect 2915 2150 2945 2202
rect 2945 2150 2957 2202
rect 2957 2150 2971 2202
rect 2995 2150 3009 2202
rect 3009 2150 3021 2202
rect 3021 2150 3051 2202
rect 3075 2150 3085 2202
rect 3085 2150 3131 2202
rect 2835 2148 2891 2150
rect 2915 2148 2971 2150
rect 2995 2148 3051 2150
rect 3075 2148 3131 2150
rect 5273 2202 5329 2204
rect 5353 2202 5409 2204
rect 5433 2202 5489 2204
rect 5513 2202 5569 2204
rect 5273 2150 5319 2202
rect 5319 2150 5329 2202
rect 5353 2150 5383 2202
rect 5383 2150 5395 2202
rect 5395 2150 5409 2202
rect 5433 2150 5447 2202
rect 5447 2150 5459 2202
rect 5459 2150 5489 2202
rect 5513 2150 5523 2202
rect 5523 2150 5569 2202
rect 5273 2148 5329 2150
rect 5353 2148 5409 2150
rect 5433 2148 5489 2150
rect 5513 2148 5569 2150
rect 7711 2202 7767 2204
rect 7791 2202 7847 2204
rect 7871 2202 7927 2204
rect 7951 2202 8007 2204
rect 7711 2150 7757 2202
rect 7757 2150 7767 2202
rect 7791 2150 7821 2202
rect 7821 2150 7833 2202
rect 7833 2150 7847 2202
rect 7871 2150 7885 2202
rect 7885 2150 7897 2202
rect 7897 2150 7927 2202
rect 7951 2150 7961 2202
rect 7961 2150 8007 2202
rect 7711 2148 7767 2150
rect 7791 2148 7847 2150
rect 7871 2148 7927 2150
rect 7951 2148 8007 2150
rect 10149 2202 10205 2204
rect 10229 2202 10285 2204
rect 10309 2202 10365 2204
rect 10389 2202 10445 2204
rect 10149 2150 10195 2202
rect 10195 2150 10205 2202
rect 10229 2150 10259 2202
rect 10259 2150 10271 2202
rect 10271 2150 10285 2202
rect 10309 2150 10323 2202
rect 10323 2150 10335 2202
rect 10335 2150 10365 2202
rect 10389 2150 10399 2202
rect 10399 2150 10445 2202
rect 10149 2148 10205 2150
rect 10229 2148 10285 2150
rect 10309 2148 10365 2150
rect 10389 2148 10445 2150
rect 9586 1128 9642 1184
rect 1766 584 1822 640
<< metal3 >>
rect 0 15330 800 15360
rect 3601 15330 3667 15333
rect 0 15328 3667 15330
rect 0 15272 3606 15328
rect 3662 15272 3667 15328
rect 0 15270 3667 15272
rect 0 15240 800 15270
rect 3601 15267 3667 15270
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 10409 14514 10475 14517
rect 11200 14514 12000 14544
rect 10409 14512 12000 14514
rect 10409 14456 10414 14512
rect 10470 14456 12000 14512
rect 10409 14454 12000 14456
rect 10409 14451 10475 14454
rect 11200 14424 12000 14454
rect 0 13698 800 13728
rect 0 13638 1594 13698
rect 0 13608 800 13638
rect 1534 13426 1594 13638
rect 2165 13632 2481 13633
rect 2165 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2481 13632
rect 2165 13567 2481 13568
rect 4603 13632 4919 13633
rect 4603 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4919 13632
rect 4603 13567 4919 13568
rect 7041 13632 7357 13633
rect 7041 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7357 13632
rect 7041 13567 7357 13568
rect 9479 13632 9795 13633
rect 9479 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9795 13632
rect 9479 13567 9795 13568
rect 3049 13426 3115 13429
rect 1534 13424 3115 13426
rect 1534 13368 3054 13424
rect 3110 13368 3115 13424
rect 1534 13366 3115 13368
rect 3049 13363 3115 13366
rect 2825 13088 3141 13089
rect 2825 13024 2831 13088
rect 2895 13024 2911 13088
rect 2975 13024 2991 13088
rect 3055 13024 3071 13088
rect 3135 13024 3141 13088
rect 2825 13023 3141 13024
rect 5263 13088 5579 13089
rect 5263 13024 5269 13088
rect 5333 13024 5349 13088
rect 5413 13024 5429 13088
rect 5493 13024 5509 13088
rect 5573 13024 5579 13088
rect 5263 13023 5579 13024
rect 7701 13088 8017 13089
rect 7701 13024 7707 13088
rect 7771 13024 7787 13088
rect 7851 13024 7867 13088
rect 7931 13024 7947 13088
rect 8011 13024 8017 13088
rect 7701 13023 8017 13024
rect 10139 13088 10455 13089
rect 10139 13024 10145 13088
rect 10209 13024 10225 13088
rect 10289 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10455 13088
rect 10139 13023 10455 13024
rect 0 12882 800 12912
rect 2681 12882 2747 12885
rect 0 12880 2747 12882
rect 0 12824 2686 12880
rect 2742 12824 2747 12880
rect 0 12822 2747 12824
rect 0 12792 800 12822
rect 2681 12819 2747 12822
rect 10409 12610 10475 12613
rect 11200 12610 12000 12640
rect 10409 12608 12000 12610
rect 10409 12552 10414 12608
rect 10470 12552 12000 12608
rect 10409 12550 12000 12552
rect 10409 12547 10475 12550
rect 2165 12544 2481 12545
rect 2165 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2481 12544
rect 2165 12479 2481 12480
rect 4603 12544 4919 12545
rect 4603 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4919 12544
rect 4603 12479 4919 12480
rect 7041 12544 7357 12545
rect 7041 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7357 12544
rect 7041 12479 7357 12480
rect 9479 12544 9795 12545
rect 9479 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9795 12544
rect 11200 12520 12000 12550
rect 9479 12479 9795 12480
rect 6085 12338 6151 12341
rect 10225 12338 10291 12341
rect 6085 12336 10291 12338
rect 6085 12280 6090 12336
rect 6146 12280 10230 12336
rect 10286 12280 10291 12336
rect 6085 12278 10291 12280
rect 6085 12275 6151 12278
rect 10225 12275 10291 12278
rect 3325 12202 3391 12205
rect 5625 12202 5691 12205
rect 6453 12202 6519 12205
rect 7097 12202 7163 12205
rect 7925 12202 7991 12205
rect 3325 12200 7163 12202
rect 3325 12144 3330 12200
rect 3386 12144 5630 12200
rect 5686 12144 6458 12200
rect 6514 12144 7102 12200
rect 7158 12144 7163 12200
rect 3325 12142 7163 12144
rect 3325 12139 3391 12142
rect 5625 12139 5691 12142
rect 6453 12139 6519 12142
rect 7097 12139 7163 12142
rect 7422 12200 7991 12202
rect 7422 12144 7930 12200
rect 7986 12144 7991 12200
rect 7422 12142 7991 12144
rect 0 12066 800 12096
rect 1669 12066 1735 12069
rect 0 12064 1735 12066
rect 0 12008 1674 12064
rect 1730 12008 1735 12064
rect 0 12006 1735 12008
rect 0 11976 800 12006
rect 1669 12003 1735 12006
rect 5717 12066 5783 12069
rect 7281 12066 7347 12069
rect 5717 12064 7347 12066
rect 5717 12008 5722 12064
rect 5778 12008 7286 12064
rect 7342 12008 7347 12064
rect 5717 12006 7347 12008
rect 5717 12003 5783 12006
rect 7281 12003 7347 12006
rect 2825 12000 3141 12001
rect 2825 11936 2831 12000
rect 2895 11936 2911 12000
rect 2975 11936 2991 12000
rect 3055 11936 3071 12000
rect 3135 11936 3141 12000
rect 2825 11935 3141 11936
rect 5263 12000 5579 12001
rect 5263 11936 5269 12000
rect 5333 11936 5349 12000
rect 5413 11936 5429 12000
rect 5493 11936 5509 12000
rect 5573 11936 5579 12000
rect 5263 11935 5579 11936
rect 7005 11930 7071 11933
rect 7422 11930 7482 12142
rect 7925 12139 7991 12142
rect 7701 12000 8017 12001
rect 7701 11936 7707 12000
rect 7771 11936 7787 12000
rect 7851 11936 7867 12000
rect 7931 11936 7947 12000
rect 8011 11936 8017 12000
rect 7701 11935 8017 11936
rect 10139 12000 10455 12001
rect 10139 11936 10145 12000
rect 10209 11936 10225 12000
rect 10289 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10455 12000
rect 10139 11935 10455 11936
rect 7005 11928 7482 11930
rect 7005 11872 7010 11928
rect 7066 11872 7482 11928
rect 7005 11870 7482 11872
rect 7005 11867 7071 11870
rect 4521 11794 4587 11797
rect 4981 11794 5047 11797
rect 4521 11792 5047 11794
rect 4521 11736 4526 11792
rect 4582 11736 4986 11792
rect 5042 11736 5047 11792
rect 4521 11734 5047 11736
rect 4521 11731 4587 11734
rect 4981 11731 5047 11734
rect 5809 11794 5875 11797
rect 6085 11794 6151 11797
rect 7373 11794 7439 11797
rect 5809 11792 7439 11794
rect 5809 11736 5814 11792
rect 5870 11736 6090 11792
rect 6146 11736 7378 11792
rect 7434 11736 7439 11792
rect 5809 11734 7439 11736
rect 5809 11731 5875 11734
rect 6085 11731 6151 11734
rect 7373 11731 7439 11734
rect 5901 11658 5967 11661
rect 7557 11658 7623 11661
rect 8201 11658 8267 11661
rect 5901 11656 8267 11658
rect 5901 11600 5906 11656
rect 5962 11600 7562 11656
rect 7618 11600 8206 11656
rect 8262 11600 8267 11656
rect 5901 11598 8267 11600
rect 5901 11595 5967 11598
rect 7557 11595 7623 11598
rect 8201 11595 8267 11598
rect 2165 11456 2481 11457
rect 2165 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2481 11456
rect 2165 11391 2481 11392
rect 4603 11456 4919 11457
rect 4603 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4919 11456
rect 4603 11391 4919 11392
rect 7041 11456 7357 11457
rect 7041 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7357 11456
rect 7041 11391 7357 11392
rect 9479 11456 9795 11457
rect 9479 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9795 11456
rect 9479 11391 9795 11392
rect 0 11250 800 11280
rect 6453 11250 6519 11253
rect 9121 11250 9187 11253
rect 0 11160 858 11250
rect 6453 11248 9187 11250
rect 6453 11192 6458 11248
rect 6514 11192 9126 11248
rect 9182 11192 9187 11248
rect 6453 11190 9187 11192
rect 6453 11187 6519 11190
rect 9121 11187 9187 11190
rect 798 11117 858 11160
rect 798 11112 907 11117
rect 798 11056 846 11112
rect 902 11056 907 11112
rect 798 11054 907 11056
rect 841 11051 907 11054
rect 2825 10912 3141 10913
rect 2825 10848 2831 10912
rect 2895 10848 2911 10912
rect 2975 10848 2991 10912
rect 3055 10848 3071 10912
rect 3135 10848 3141 10912
rect 2825 10847 3141 10848
rect 5263 10912 5579 10913
rect 5263 10848 5269 10912
rect 5333 10848 5349 10912
rect 5413 10848 5429 10912
rect 5493 10848 5509 10912
rect 5573 10848 5579 10912
rect 5263 10847 5579 10848
rect 7701 10912 8017 10913
rect 7701 10848 7707 10912
rect 7771 10848 7787 10912
rect 7851 10848 7867 10912
rect 7931 10848 7947 10912
rect 8011 10848 8017 10912
rect 7701 10847 8017 10848
rect 10139 10912 10455 10913
rect 10139 10848 10145 10912
rect 10209 10848 10225 10912
rect 10289 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10455 10912
rect 10139 10847 10455 10848
rect 3969 10706 4035 10709
rect 4429 10706 4495 10709
rect 5441 10706 5507 10709
rect 3969 10704 5507 10706
rect 3969 10648 3974 10704
rect 4030 10648 4434 10704
rect 4490 10648 5446 10704
rect 5502 10648 5507 10704
rect 3969 10646 5507 10648
rect 3969 10643 4035 10646
rect 4429 10643 4495 10646
rect 5441 10643 5507 10646
rect 10409 10706 10475 10709
rect 11200 10706 12000 10736
rect 10409 10704 12000 10706
rect 10409 10648 10414 10704
rect 10470 10648 12000 10704
rect 10409 10646 12000 10648
rect 10409 10643 10475 10646
rect 11200 10616 12000 10646
rect 841 10570 907 10573
rect 798 10568 907 10570
rect 798 10512 846 10568
rect 902 10512 907 10568
rect 798 10507 907 10512
rect 798 10464 858 10507
rect 0 10374 858 10464
rect 0 10344 800 10374
rect 2165 10368 2481 10369
rect 2165 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2481 10368
rect 2165 10303 2481 10304
rect 4603 10368 4919 10369
rect 4603 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4919 10368
rect 4603 10303 4919 10304
rect 7041 10368 7357 10369
rect 7041 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7357 10368
rect 7041 10303 7357 10304
rect 9479 10368 9795 10369
rect 9479 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9795 10368
rect 9479 10303 9795 10304
rect 2825 9824 3141 9825
rect 2825 9760 2831 9824
rect 2895 9760 2911 9824
rect 2975 9760 2991 9824
rect 3055 9760 3071 9824
rect 3135 9760 3141 9824
rect 2825 9759 3141 9760
rect 5263 9824 5579 9825
rect 5263 9760 5269 9824
rect 5333 9760 5349 9824
rect 5413 9760 5429 9824
rect 5493 9760 5509 9824
rect 5573 9760 5579 9824
rect 5263 9759 5579 9760
rect 7701 9824 8017 9825
rect 7701 9760 7707 9824
rect 7771 9760 7787 9824
rect 7851 9760 7867 9824
rect 7931 9760 7947 9824
rect 8011 9760 8017 9824
rect 7701 9759 8017 9760
rect 10139 9824 10455 9825
rect 10139 9760 10145 9824
rect 10209 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10455 9824
rect 10139 9759 10455 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 841 8938 907 8941
rect 798 8936 907 8938
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8875 907 8880
rect 5717 8938 5783 8941
rect 6177 8938 6243 8941
rect 5717 8936 6243 8938
rect 5717 8880 5722 8936
rect 5778 8880 6182 8936
rect 6238 8880 6243 8936
rect 5717 8878 6243 8880
rect 5717 8875 5783 8878
rect 6177 8875 6243 8878
rect 798 8832 858 8875
rect 0 8742 858 8832
rect 10869 8802 10935 8805
rect 11200 8802 12000 8832
rect 10869 8800 12000 8802
rect 10869 8744 10874 8800
rect 10930 8744 12000 8800
rect 10869 8742 12000 8744
rect 0 8712 800 8742
rect 10869 8739 10935 8742
rect 2825 8736 3141 8737
rect 2825 8672 2831 8736
rect 2895 8672 2911 8736
rect 2975 8672 2991 8736
rect 3055 8672 3071 8736
rect 3135 8672 3141 8736
rect 2825 8671 3141 8672
rect 5263 8736 5579 8737
rect 5263 8672 5269 8736
rect 5333 8672 5349 8736
rect 5413 8672 5429 8736
rect 5493 8672 5509 8736
rect 5573 8672 5579 8736
rect 5263 8671 5579 8672
rect 7701 8736 8017 8737
rect 7701 8672 7707 8736
rect 7771 8672 7787 8736
rect 7851 8672 7867 8736
rect 7931 8672 7947 8736
rect 8011 8672 8017 8736
rect 7701 8671 8017 8672
rect 10139 8736 10455 8737
rect 10139 8672 10145 8736
rect 10209 8672 10225 8736
rect 10289 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10455 8736
rect 11200 8712 12000 8742
rect 10139 8671 10455 8672
rect 5993 8394 6059 8397
rect 6269 8394 6335 8397
rect 8385 8394 8451 8397
rect 5993 8392 8451 8394
rect 5993 8336 5998 8392
rect 6054 8336 6274 8392
rect 6330 8336 8390 8392
rect 8446 8336 8451 8392
rect 5993 8334 8451 8336
rect 5993 8331 6059 8334
rect 6269 8331 6335 8334
rect 8385 8331 8451 8334
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7986 800 8016
rect 1393 7986 1459 7989
rect 0 7984 1459 7986
rect 0 7928 1398 7984
rect 1454 7928 1459 7984
rect 0 7926 1459 7928
rect 0 7896 800 7926
rect 1393 7923 1459 7926
rect 2825 7648 3141 7649
rect 2825 7584 2831 7648
rect 2895 7584 2911 7648
rect 2975 7584 2991 7648
rect 3055 7584 3071 7648
rect 3135 7584 3141 7648
rect 2825 7583 3141 7584
rect 5263 7648 5579 7649
rect 5263 7584 5269 7648
rect 5333 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5579 7648
rect 5263 7583 5579 7584
rect 7701 7648 8017 7649
rect 7701 7584 7707 7648
rect 7771 7584 7787 7648
rect 7851 7584 7867 7648
rect 7931 7584 7947 7648
rect 8011 7584 8017 7648
rect 7701 7583 8017 7584
rect 10139 7648 10455 7649
rect 10139 7584 10145 7648
rect 10209 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10455 7648
rect 10139 7583 10455 7584
rect 6085 7442 6151 7445
rect 2730 7440 6151 7442
rect 2730 7384 6090 7440
rect 6146 7384 6151 7440
rect 2730 7382 6151 7384
rect 841 7306 907 7309
rect 798 7304 907 7306
rect 798 7248 846 7304
rect 902 7248 907 7304
rect 798 7243 907 7248
rect 1577 7306 1643 7309
rect 2730 7306 2790 7382
rect 6085 7379 6151 7382
rect 1577 7304 2790 7306
rect 1577 7248 1582 7304
rect 1638 7248 2790 7304
rect 1577 7246 2790 7248
rect 1577 7243 1643 7246
rect 798 7200 858 7243
rect 0 7110 858 7200
rect 0 7080 800 7110
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 2957 6898 3023 6901
rect 3509 6898 3575 6901
rect 5901 6898 5967 6901
rect 2957 6896 5967 6898
rect 2957 6840 2962 6896
rect 3018 6840 3514 6896
rect 3570 6840 5906 6896
rect 5962 6840 5967 6896
rect 2957 6838 5967 6840
rect 2957 6835 3023 6838
rect 3509 6835 3575 6838
rect 5901 6835 5967 6838
rect 10409 6898 10475 6901
rect 11200 6898 12000 6928
rect 10409 6896 12000 6898
rect 10409 6840 10414 6896
rect 10470 6840 12000 6896
rect 10409 6838 12000 6840
rect 10409 6835 10475 6838
rect 11200 6808 12000 6838
rect 5257 6762 5323 6765
rect 5809 6762 5875 6765
rect 6269 6762 6335 6765
rect 5257 6760 6335 6762
rect 5257 6704 5262 6760
rect 5318 6704 5814 6760
rect 5870 6704 6274 6760
rect 6330 6704 6335 6760
rect 5257 6702 6335 6704
rect 5257 6699 5323 6702
rect 5809 6699 5875 6702
rect 6269 6699 6335 6702
rect 2825 6560 3141 6561
rect 2825 6496 2831 6560
rect 2895 6496 2911 6560
rect 2975 6496 2991 6560
rect 3055 6496 3071 6560
rect 3135 6496 3141 6560
rect 2825 6495 3141 6496
rect 5263 6560 5579 6561
rect 5263 6496 5269 6560
rect 5333 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5579 6560
rect 5263 6495 5579 6496
rect 7701 6560 8017 6561
rect 7701 6496 7707 6560
rect 7771 6496 7787 6560
rect 7851 6496 7867 6560
rect 7931 6496 7947 6560
rect 8011 6496 8017 6560
rect 7701 6495 8017 6496
rect 10139 6560 10455 6561
rect 10139 6496 10145 6560
rect 10209 6496 10225 6560
rect 10289 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10455 6560
rect 10139 6495 10455 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 0 6264 800 6294
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 2825 5472 3141 5473
rect 2825 5408 2831 5472
rect 2895 5408 2911 5472
rect 2975 5408 2991 5472
rect 3055 5408 3071 5472
rect 3135 5408 3141 5472
rect 2825 5407 3141 5408
rect 5263 5472 5579 5473
rect 5263 5408 5269 5472
rect 5333 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5579 5472
rect 5263 5407 5579 5408
rect 7701 5472 8017 5473
rect 7701 5408 7707 5472
rect 7771 5408 7787 5472
rect 7851 5408 7867 5472
rect 7931 5408 7947 5472
rect 8011 5408 8017 5472
rect 7701 5407 8017 5408
rect 10139 5472 10455 5473
rect 10139 5408 10145 5472
rect 10209 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10455 5472
rect 10139 5407 10455 5408
rect 10409 4994 10475 4997
rect 11200 4994 12000 5024
rect 10409 4992 12000 4994
rect 10409 4936 10414 4992
rect 10470 4936 12000 4992
rect 10409 4934 12000 4936
rect 10409 4931 10475 4934
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 11200 4904 12000 4934
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 0 4632 858 4722
rect 798 4589 858 4632
rect 798 4584 907 4589
rect 798 4528 846 4584
rect 902 4528 907 4584
rect 798 4526 907 4528
rect 841 4523 907 4526
rect 2825 4384 3141 4385
rect 2825 4320 2831 4384
rect 2895 4320 2911 4384
rect 2975 4320 2991 4384
rect 3055 4320 3071 4384
rect 3135 4320 3141 4384
rect 2825 4319 3141 4320
rect 5263 4384 5579 4385
rect 5263 4320 5269 4384
rect 5333 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5579 4384
rect 5263 4319 5579 4320
rect 7701 4384 8017 4385
rect 7701 4320 7707 4384
rect 7771 4320 7787 4384
rect 7851 4320 7867 4384
rect 7931 4320 7947 4384
rect 8011 4320 8017 4384
rect 7701 4319 8017 4320
rect 10139 4384 10455 4385
rect 10139 4320 10145 4384
rect 10209 4320 10225 4384
rect 10289 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10455 4384
rect 10139 4319 10455 4320
rect 2313 4178 2379 4181
rect 6913 4178 6979 4181
rect 2313 4176 6979 4178
rect 2313 4120 2318 4176
rect 2374 4120 6918 4176
rect 6974 4120 6979 4176
rect 2313 4118 6979 4120
rect 2313 4115 2379 4118
rect 6913 4115 6979 4118
rect 841 4042 907 4045
rect 798 4040 907 4042
rect 798 3984 846 4040
rect 902 3984 907 4040
rect 798 3979 907 3984
rect 798 3936 858 3979
rect 0 3846 858 3936
rect 0 3816 800 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 4705 3634 4771 3637
rect 6177 3634 6243 3637
rect 4705 3632 6243 3634
rect 4705 3576 4710 3632
rect 4766 3576 6182 3632
rect 6238 3576 6243 3632
rect 4705 3574 6243 3576
rect 4705 3571 4771 3574
rect 6177 3571 6243 3574
rect 3877 3498 3943 3501
rect 9213 3498 9279 3501
rect 3877 3496 9279 3498
rect 3877 3440 3882 3496
rect 3938 3440 9218 3496
rect 9274 3440 9279 3496
rect 3877 3438 9279 3440
rect 3877 3435 3943 3438
rect 9213 3435 9279 3438
rect 2825 3296 3141 3297
rect 2825 3232 2831 3296
rect 2895 3232 2911 3296
rect 2975 3232 2991 3296
rect 3055 3232 3071 3296
rect 3135 3232 3141 3296
rect 2825 3231 3141 3232
rect 5263 3296 5579 3297
rect 5263 3232 5269 3296
rect 5333 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5579 3296
rect 5263 3231 5579 3232
rect 7701 3296 8017 3297
rect 7701 3232 7707 3296
rect 7771 3232 7787 3296
rect 7851 3232 7867 3296
rect 7931 3232 7947 3296
rect 8011 3232 8017 3296
rect 7701 3231 8017 3232
rect 10139 3296 10455 3297
rect 10139 3232 10145 3296
rect 10209 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10455 3296
rect 10139 3231 10455 3232
rect 841 3226 907 3229
rect 798 3224 907 3226
rect 798 3168 846 3224
rect 902 3168 907 3224
rect 798 3163 907 3168
rect 798 3120 858 3163
rect 0 3030 858 3120
rect 1945 3090 2011 3093
rect 6361 3090 6427 3093
rect 1945 3088 6427 3090
rect 1945 3032 1950 3088
rect 2006 3032 6366 3088
rect 6422 3032 6427 3088
rect 1945 3030 6427 3032
rect 0 3000 800 3030
rect 1945 3027 2011 3030
rect 6361 3027 6427 3030
rect 6637 3090 6703 3093
rect 7741 3090 7807 3093
rect 6637 3088 7807 3090
rect 6637 3032 6642 3088
rect 6698 3032 7746 3088
rect 7802 3032 7807 3088
rect 6637 3030 7807 3032
rect 6637 3027 6703 3030
rect 7741 3027 7807 3030
rect 10501 3090 10567 3093
rect 11200 3090 12000 3120
rect 10501 3088 12000 3090
rect 10501 3032 10506 3088
rect 10562 3032 12000 3088
rect 10501 3030 12000 3032
rect 10501 3027 10567 3030
rect 11200 3000 12000 3030
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 0 2184 800 2214
rect 2825 2208 3141 2209
rect 2825 2144 2831 2208
rect 2895 2144 2911 2208
rect 2975 2144 2991 2208
rect 3055 2144 3071 2208
rect 3135 2144 3141 2208
rect 2825 2143 3141 2144
rect 5263 2208 5579 2209
rect 5263 2144 5269 2208
rect 5333 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5579 2208
rect 5263 2143 5579 2144
rect 7701 2208 8017 2209
rect 7701 2144 7707 2208
rect 7771 2144 7787 2208
rect 7851 2144 7867 2208
rect 7931 2144 7947 2208
rect 8011 2144 8017 2208
rect 7701 2143 8017 2144
rect 10139 2208 10455 2209
rect 10139 2144 10145 2208
rect 10209 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10455 2208
rect 10139 2143 10455 2144
rect 0 1458 800 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 800 1398
rect 1485 1395 1551 1398
rect 9581 1186 9647 1189
rect 11200 1186 12000 1216
rect 9581 1184 12000 1186
rect 9581 1128 9586 1184
rect 9642 1128 12000 1184
rect 9581 1126 12000 1128
rect 9581 1123 9647 1126
rect 11200 1096 12000 1126
rect 0 642 800 672
rect 1761 642 1827 645
rect 0 640 1827 642
rect 0 584 1766 640
rect 1822 584 1827 640
rect 0 582 1827 584
rect 0 552 800 582
rect 1761 579 1827 582
<< via3 >>
rect 2171 13628 2235 13632
rect 2171 13572 2175 13628
rect 2175 13572 2231 13628
rect 2231 13572 2235 13628
rect 2171 13568 2235 13572
rect 2251 13628 2315 13632
rect 2251 13572 2255 13628
rect 2255 13572 2311 13628
rect 2311 13572 2315 13628
rect 2251 13568 2315 13572
rect 2331 13628 2395 13632
rect 2331 13572 2335 13628
rect 2335 13572 2391 13628
rect 2391 13572 2395 13628
rect 2331 13568 2395 13572
rect 2411 13628 2475 13632
rect 2411 13572 2415 13628
rect 2415 13572 2471 13628
rect 2471 13572 2475 13628
rect 2411 13568 2475 13572
rect 4609 13628 4673 13632
rect 4609 13572 4613 13628
rect 4613 13572 4669 13628
rect 4669 13572 4673 13628
rect 4609 13568 4673 13572
rect 4689 13628 4753 13632
rect 4689 13572 4693 13628
rect 4693 13572 4749 13628
rect 4749 13572 4753 13628
rect 4689 13568 4753 13572
rect 4769 13628 4833 13632
rect 4769 13572 4773 13628
rect 4773 13572 4829 13628
rect 4829 13572 4833 13628
rect 4769 13568 4833 13572
rect 4849 13628 4913 13632
rect 4849 13572 4853 13628
rect 4853 13572 4909 13628
rect 4909 13572 4913 13628
rect 4849 13568 4913 13572
rect 7047 13628 7111 13632
rect 7047 13572 7051 13628
rect 7051 13572 7107 13628
rect 7107 13572 7111 13628
rect 7047 13568 7111 13572
rect 7127 13628 7191 13632
rect 7127 13572 7131 13628
rect 7131 13572 7187 13628
rect 7187 13572 7191 13628
rect 7127 13568 7191 13572
rect 7207 13628 7271 13632
rect 7207 13572 7211 13628
rect 7211 13572 7267 13628
rect 7267 13572 7271 13628
rect 7207 13568 7271 13572
rect 7287 13628 7351 13632
rect 7287 13572 7291 13628
rect 7291 13572 7347 13628
rect 7347 13572 7351 13628
rect 7287 13568 7351 13572
rect 9485 13628 9549 13632
rect 9485 13572 9489 13628
rect 9489 13572 9545 13628
rect 9545 13572 9549 13628
rect 9485 13568 9549 13572
rect 9565 13628 9629 13632
rect 9565 13572 9569 13628
rect 9569 13572 9625 13628
rect 9625 13572 9629 13628
rect 9565 13568 9629 13572
rect 9645 13628 9709 13632
rect 9645 13572 9649 13628
rect 9649 13572 9705 13628
rect 9705 13572 9709 13628
rect 9645 13568 9709 13572
rect 9725 13628 9789 13632
rect 9725 13572 9729 13628
rect 9729 13572 9785 13628
rect 9785 13572 9789 13628
rect 9725 13568 9789 13572
rect 2831 13084 2895 13088
rect 2831 13028 2835 13084
rect 2835 13028 2891 13084
rect 2891 13028 2895 13084
rect 2831 13024 2895 13028
rect 2911 13084 2975 13088
rect 2911 13028 2915 13084
rect 2915 13028 2971 13084
rect 2971 13028 2975 13084
rect 2911 13024 2975 13028
rect 2991 13084 3055 13088
rect 2991 13028 2995 13084
rect 2995 13028 3051 13084
rect 3051 13028 3055 13084
rect 2991 13024 3055 13028
rect 3071 13084 3135 13088
rect 3071 13028 3075 13084
rect 3075 13028 3131 13084
rect 3131 13028 3135 13084
rect 3071 13024 3135 13028
rect 5269 13084 5333 13088
rect 5269 13028 5273 13084
rect 5273 13028 5329 13084
rect 5329 13028 5333 13084
rect 5269 13024 5333 13028
rect 5349 13084 5413 13088
rect 5349 13028 5353 13084
rect 5353 13028 5409 13084
rect 5409 13028 5413 13084
rect 5349 13024 5413 13028
rect 5429 13084 5493 13088
rect 5429 13028 5433 13084
rect 5433 13028 5489 13084
rect 5489 13028 5493 13084
rect 5429 13024 5493 13028
rect 5509 13084 5573 13088
rect 5509 13028 5513 13084
rect 5513 13028 5569 13084
rect 5569 13028 5573 13084
rect 5509 13024 5573 13028
rect 7707 13084 7771 13088
rect 7707 13028 7711 13084
rect 7711 13028 7767 13084
rect 7767 13028 7771 13084
rect 7707 13024 7771 13028
rect 7787 13084 7851 13088
rect 7787 13028 7791 13084
rect 7791 13028 7847 13084
rect 7847 13028 7851 13084
rect 7787 13024 7851 13028
rect 7867 13084 7931 13088
rect 7867 13028 7871 13084
rect 7871 13028 7927 13084
rect 7927 13028 7931 13084
rect 7867 13024 7931 13028
rect 7947 13084 8011 13088
rect 7947 13028 7951 13084
rect 7951 13028 8007 13084
rect 8007 13028 8011 13084
rect 7947 13024 8011 13028
rect 10145 13084 10209 13088
rect 10145 13028 10149 13084
rect 10149 13028 10205 13084
rect 10205 13028 10209 13084
rect 10145 13024 10209 13028
rect 10225 13084 10289 13088
rect 10225 13028 10229 13084
rect 10229 13028 10285 13084
rect 10285 13028 10289 13084
rect 10225 13024 10289 13028
rect 10305 13084 10369 13088
rect 10305 13028 10309 13084
rect 10309 13028 10365 13084
rect 10365 13028 10369 13084
rect 10305 13024 10369 13028
rect 10385 13084 10449 13088
rect 10385 13028 10389 13084
rect 10389 13028 10445 13084
rect 10445 13028 10449 13084
rect 10385 13024 10449 13028
rect 2171 12540 2235 12544
rect 2171 12484 2175 12540
rect 2175 12484 2231 12540
rect 2231 12484 2235 12540
rect 2171 12480 2235 12484
rect 2251 12540 2315 12544
rect 2251 12484 2255 12540
rect 2255 12484 2311 12540
rect 2311 12484 2315 12540
rect 2251 12480 2315 12484
rect 2331 12540 2395 12544
rect 2331 12484 2335 12540
rect 2335 12484 2391 12540
rect 2391 12484 2395 12540
rect 2331 12480 2395 12484
rect 2411 12540 2475 12544
rect 2411 12484 2415 12540
rect 2415 12484 2471 12540
rect 2471 12484 2475 12540
rect 2411 12480 2475 12484
rect 4609 12540 4673 12544
rect 4609 12484 4613 12540
rect 4613 12484 4669 12540
rect 4669 12484 4673 12540
rect 4609 12480 4673 12484
rect 4689 12540 4753 12544
rect 4689 12484 4693 12540
rect 4693 12484 4749 12540
rect 4749 12484 4753 12540
rect 4689 12480 4753 12484
rect 4769 12540 4833 12544
rect 4769 12484 4773 12540
rect 4773 12484 4829 12540
rect 4829 12484 4833 12540
rect 4769 12480 4833 12484
rect 4849 12540 4913 12544
rect 4849 12484 4853 12540
rect 4853 12484 4909 12540
rect 4909 12484 4913 12540
rect 4849 12480 4913 12484
rect 7047 12540 7111 12544
rect 7047 12484 7051 12540
rect 7051 12484 7107 12540
rect 7107 12484 7111 12540
rect 7047 12480 7111 12484
rect 7127 12540 7191 12544
rect 7127 12484 7131 12540
rect 7131 12484 7187 12540
rect 7187 12484 7191 12540
rect 7127 12480 7191 12484
rect 7207 12540 7271 12544
rect 7207 12484 7211 12540
rect 7211 12484 7267 12540
rect 7267 12484 7271 12540
rect 7207 12480 7271 12484
rect 7287 12540 7351 12544
rect 7287 12484 7291 12540
rect 7291 12484 7347 12540
rect 7347 12484 7351 12540
rect 7287 12480 7351 12484
rect 9485 12540 9549 12544
rect 9485 12484 9489 12540
rect 9489 12484 9545 12540
rect 9545 12484 9549 12540
rect 9485 12480 9549 12484
rect 9565 12540 9629 12544
rect 9565 12484 9569 12540
rect 9569 12484 9625 12540
rect 9625 12484 9629 12540
rect 9565 12480 9629 12484
rect 9645 12540 9709 12544
rect 9645 12484 9649 12540
rect 9649 12484 9705 12540
rect 9705 12484 9709 12540
rect 9645 12480 9709 12484
rect 9725 12540 9789 12544
rect 9725 12484 9729 12540
rect 9729 12484 9785 12540
rect 9785 12484 9789 12540
rect 9725 12480 9789 12484
rect 2831 11996 2895 12000
rect 2831 11940 2835 11996
rect 2835 11940 2891 11996
rect 2891 11940 2895 11996
rect 2831 11936 2895 11940
rect 2911 11996 2975 12000
rect 2911 11940 2915 11996
rect 2915 11940 2971 11996
rect 2971 11940 2975 11996
rect 2911 11936 2975 11940
rect 2991 11996 3055 12000
rect 2991 11940 2995 11996
rect 2995 11940 3051 11996
rect 3051 11940 3055 11996
rect 2991 11936 3055 11940
rect 3071 11996 3135 12000
rect 3071 11940 3075 11996
rect 3075 11940 3131 11996
rect 3131 11940 3135 11996
rect 3071 11936 3135 11940
rect 5269 11996 5333 12000
rect 5269 11940 5273 11996
rect 5273 11940 5329 11996
rect 5329 11940 5333 11996
rect 5269 11936 5333 11940
rect 5349 11996 5413 12000
rect 5349 11940 5353 11996
rect 5353 11940 5409 11996
rect 5409 11940 5413 11996
rect 5349 11936 5413 11940
rect 5429 11996 5493 12000
rect 5429 11940 5433 11996
rect 5433 11940 5489 11996
rect 5489 11940 5493 11996
rect 5429 11936 5493 11940
rect 5509 11996 5573 12000
rect 5509 11940 5513 11996
rect 5513 11940 5569 11996
rect 5569 11940 5573 11996
rect 5509 11936 5573 11940
rect 7707 11996 7771 12000
rect 7707 11940 7711 11996
rect 7711 11940 7767 11996
rect 7767 11940 7771 11996
rect 7707 11936 7771 11940
rect 7787 11996 7851 12000
rect 7787 11940 7791 11996
rect 7791 11940 7847 11996
rect 7847 11940 7851 11996
rect 7787 11936 7851 11940
rect 7867 11996 7931 12000
rect 7867 11940 7871 11996
rect 7871 11940 7927 11996
rect 7927 11940 7931 11996
rect 7867 11936 7931 11940
rect 7947 11996 8011 12000
rect 7947 11940 7951 11996
rect 7951 11940 8007 11996
rect 8007 11940 8011 11996
rect 7947 11936 8011 11940
rect 10145 11996 10209 12000
rect 10145 11940 10149 11996
rect 10149 11940 10205 11996
rect 10205 11940 10209 11996
rect 10145 11936 10209 11940
rect 10225 11996 10289 12000
rect 10225 11940 10229 11996
rect 10229 11940 10285 11996
rect 10285 11940 10289 11996
rect 10225 11936 10289 11940
rect 10305 11996 10369 12000
rect 10305 11940 10309 11996
rect 10309 11940 10365 11996
rect 10365 11940 10369 11996
rect 10305 11936 10369 11940
rect 10385 11996 10449 12000
rect 10385 11940 10389 11996
rect 10389 11940 10445 11996
rect 10445 11940 10449 11996
rect 10385 11936 10449 11940
rect 2171 11452 2235 11456
rect 2171 11396 2175 11452
rect 2175 11396 2231 11452
rect 2231 11396 2235 11452
rect 2171 11392 2235 11396
rect 2251 11452 2315 11456
rect 2251 11396 2255 11452
rect 2255 11396 2311 11452
rect 2311 11396 2315 11452
rect 2251 11392 2315 11396
rect 2331 11452 2395 11456
rect 2331 11396 2335 11452
rect 2335 11396 2391 11452
rect 2391 11396 2395 11452
rect 2331 11392 2395 11396
rect 2411 11452 2475 11456
rect 2411 11396 2415 11452
rect 2415 11396 2471 11452
rect 2471 11396 2475 11452
rect 2411 11392 2475 11396
rect 4609 11452 4673 11456
rect 4609 11396 4613 11452
rect 4613 11396 4669 11452
rect 4669 11396 4673 11452
rect 4609 11392 4673 11396
rect 4689 11452 4753 11456
rect 4689 11396 4693 11452
rect 4693 11396 4749 11452
rect 4749 11396 4753 11452
rect 4689 11392 4753 11396
rect 4769 11452 4833 11456
rect 4769 11396 4773 11452
rect 4773 11396 4829 11452
rect 4829 11396 4833 11452
rect 4769 11392 4833 11396
rect 4849 11452 4913 11456
rect 4849 11396 4853 11452
rect 4853 11396 4909 11452
rect 4909 11396 4913 11452
rect 4849 11392 4913 11396
rect 7047 11452 7111 11456
rect 7047 11396 7051 11452
rect 7051 11396 7107 11452
rect 7107 11396 7111 11452
rect 7047 11392 7111 11396
rect 7127 11452 7191 11456
rect 7127 11396 7131 11452
rect 7131 11396 7187 11452
rect 7187 11396 7191 11452
rect 7127 11392 7191 11396
rect 7207 11452 7271 11456
rect 7207 11396 7211 11452
rect 7211 11396 7267 11452
rect 7267 11396 7271 11452
rect 7207 11392 7271 11396
rect 7287 11452 7351 11456
rect 7287 11396 7291 11452
rect 7291 11396 7347 11452
rect 7347 11396 7351 11452
rect 7287 11392 7351 11396
rect 9485 11452 9549 11456
rect 9485 11396 9489 11452
rect 9489 11396 9545 11452
rect 9545 11396 9549 11452
rect 9485 11392 9549 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 2831 10908 2895 10912
rect 2831 10852 2835 10908
rect 2835 10852 2891 10908
rect 2891 10852 2895 10908
rect 2831 10848 2895 10852
rect 2911 10908 2975 10912
rect 2911 10852 2915 10908
rect 2915 10852 2971 10908
rect 2971 10852 2975 10908
rect 2911 10848 2975 10852
rect 2991 10908 3055 10912
rect 2991 10852 2995 10908
rect 2995 10852 3051 10908
rect 3051 10852 3055 10908
rect 2991 10848 3055 10852
rect 3071 10908 3135 10912
rect 3071 10852 3075 10908
rect 3075 10852 3131 10908
rect 3131 10852 3135 10908
rect 3071 10848 3135 10852
rect 5269 10908 5333 10912
rect 5269 10852 5273 10908
rect 5273 10852 5329 10908
rect 5329 10852 5333 10908
rect 5269 10848 5333 10852
rect 5349 10908 5413 10912
rect 5349 10852 5353 10908
rect 5353 10852 5409 10908
rect 5409 10852 5413 10908
rect 5349 10848 5413 10852
rect 5429 10908 5493 10912
rect 5429 10852 5433 10908
rect 5433 10852 5489 10908
rect 5489 10852 5493 10908
rect 5429 10848 5493 10852
rect 5509 10908 5573 10912
rect 5509 10852 5513 10908
rect 5513 10852 5569 10908
rect 5569 10852 5573 10908
rect 5509 10848 5573 10852
rect 7707 10908 7771 10912
rect 7707 10852 7711 10908
rect 7711 10852 7767 10908
rect 7767 10852 7771 10908
rect 7707 10848 7771 10852
rect 7787 10908 7851 10912
rect 7787 10852 7791 10908
rect 7791 10852 7847 10908
rect 7847 10852 7851 10908
rect 7787 10848 7851 10852
rect 7867 10908 7931 10912
rect 7867 10852 7871 10908
rect 7871 10852 7927 10908
rect 7927 10852 7931 10908
rect 7867 10848 7931 10852
rect 7947 10908 8011 10912
rect 7947 10852 7951 10908
rect 7951 10852 8007 10908
rect 8007 10852 8011 10908
rect 7947 10848 8011 10852
rect 10145 10908 10209 10912
rect 10145 10852 10149 10908
rect 10149 10852 10205 10908
rect 10205 10852 10209 10908
rect 10145 10848 10209 10852
rect 10225 10908 10289 10912
rect 10225 10852 10229 10908
rect 10229 10852 10285 10908
rect 10285 10852 10289 10908
rect 10225 10848 10289 10852
rect 10305 10908 10369 10912
rect 10305 10852 10309 10908
rect 10309 10852 10365 10908
rect 10365 10852 10369 10908
rect 10305 10848 10369 10852
rect 10385 10908 10449 10912
rect 10385 10852 10389 10908
rect 10389 10852 10445 10908
rect 10445 10852 10449 10908
rect 10385 10848 10449 10852
rect 2171 10364 2235 10368
rect 2171 10308 2175 10364
rect 2175 10308 2231 10364
rect 2231 10308 2235 10364
rect 2171 10304 2235 10308
rect 2251 10364 2315 10368
rect 2251 10308 2255 10364
rect 2255 10308 2311 10364
rect 2311 10308 2315 10364
rect 2251 10304 2315 10308
rect 2331 10364 2395 10368
rect 2331 10308 2335 10364
rect 2335 10308 2391 10364
rect 2391 10308 2395 10364
rect 2331 10304 2395 10308
rect 2411 10364 2475 10368
rect 2411 10308 2415 10364
rect 2415 10308 2471 10364
rect 2471 10308 2475 10364
rect 2411 10304 2475 10308
rect 4609 10364 4673 10368
rect 4609 10308 4613 10364
rect 4613 10308 4669 10364
rect 4669 10308 4673 10364
rect 4609 10304 4673 10308
rect 4689 10364 4753 10368
rect 4689 10308 4693 10364
rect 4693 10308 4749 10364
rect 4749 10308 4753 10364
rect 4689 10304 4753 10308
rect 4769 10364 4833 10368
rect 4769 10308 4773 10364
rect 4773 10308 4829 10364
rect 4829 10308 4833 10364
rect 4769 10304 4833 10308
rect 4849 10364 4913 10368
rect 4849 10308 4853 10364
rect 4853 10308 4909 10364
rect 4909 10308 4913 10364
rect 4849 10304 4913 10308
rect 7047 10364 7111 10368
rect 7047 10308 7051 10364
rect 7051 10308 7107 10364
rect 7107 10308 7111 10364
rect 7047 10304 7111 10308
rect 7127 10364 7191 10368
rect 7127 10308 7131 10364
rect 7131 10308 7187 10364
rect 7187 10308 7191 10364
rect 7127 10304 7191 10308
rect 7207 10364 7271 10368
rect 7207 10308 7211 10364
rect 7211 10308 7267 10364
rect 7267 10308 7271 10364
rect 7207 10304 7271 10308
rect 7287 10364 7351 10368
rect 7287 10308 7291 10364
rect 7291 10308 7347 10364
rect 7347 10308 7351 10364
rect 7287 10304 7351 10308
rect 9485 10364 9549 10368
rect 9485 10308 9489 10364
rect 9489 10308 9545 10364
rect 9545 10308 9549 10364
rect 9485 10304 9549 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 2831 9820 2895 9824
rect 2831 9764 2835 9820
rect 2835 9764 2891 9820
rect 2891 9764 2895 9820
rect 2831 9760 2895 9764
rect 2911 9820 2975 9824
rect 2911 9764 2915 9820
rect 2915 9764 2971 9820
rect 2971 9764 2975 9820
rect 2911 9760 2975 9764
rect 2991 9820 3055 9824
rect 2991 9764 2995 9820
rect 2995 9764 3051 9820
rect 3051 9764 3055 9820
rect 2991 9760 3055 9764
rect 3071 9820 3135 9824
rect 3071 9764 3075 9820
rect 3075 9764 3131 9820
rect 3131 9764 3135 9820
rect 3071 9760 3135 9764
rect 5269 9820 5333 9824
rect 5269 9764 5273 9820
rect 5273 9764 5329 9820
rect 5329 9764 5333 9820
rect 5269 9760 5333 9764
rect 5349 9820 5413 9824
rect 5349 9764 5353 9820
rect 5353 9764 5409 9820
rect 5409 9764 5413 9820
rect 5349 9760 5413 9764
rect 5429 9820 5493 9824
rect 5429 9764 5433 9820
rect 5433 9764 5489 9820
rect 5489 9764 5493 9820
rect 5429 9760 5493 9764
rect 5509 9820 5573 9824
rect 5509 9764 5513 9820
rect 5513 9764 5569 9820
rect 5569 9764 5573 9820
rect 5509 9760 5573 9764
rect 7707 9820 7771 9824
rect 7707 9764 7711 9820
rect 7711 9764 7767 9820
rect 7767 9764 7771 9820
rect 7707 9760 7771 9764
rect 7787 9820 7851 9824
rect 7787 9764 7791 9820
rect 7791 9764 7847 9820
rect 7847 9764 7851 9820
rect 7787 9760 7851 9764
rect 7867 9820 7931 9824
rect 7867 9764 7871 9820
rect 7871 9764 7927 9820
rect 7927 9764 7931 9820
rect 7867 9760 7931 9764
rect 7947 9820 8011 9824
rect 7947 9764 7951 9820
rect 7951 9764 8007 9820
rect 8007 9764 8011 9820
rect 7947 9760 8011 9764
rect 10145 9820 10209 9824
rect 10145 9764 10149 9820
rect 10149 9764 10205 9820
rect 10205 9764 10209 9820
rect 10145 9760 10209 9764
rect 10225 9820 10289 9824
rect 10225 9764 10229 9820
rect 10229 9764 10285 9820
rect 10285 9764 10289 9820
rect 10225 9760 10289 9764
rect 10305 9820 10369 9824
rect 10305 9764 10309 9820
rect 10309 9764 10365 9820
rect 10365 9764 10369 9820
rect 10305 9760 10369 9764
rect 10385 9820 10449 9824
rect 10385 9764 10389 9820
rect 10389 9764 10445 9820
rect 10445 9764 10449 9820
rect 10385 9760 10449 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 2831 8732 2895 8736
rect 2831 8676 2835 8732
rect 2835 8676 2891 8732
rect 2891 8676 2895 8732
rect 2831 8672 2895 8676
rect 2911 8732 2975 8736
rect 2911 8676 2915 8732
rect 2915 8676 2971 8732
rect 2971 8676 2975 8732
rect 2911 8672 2975 8676
rect 2991 8732 3055 8736
rect 2991 8676 2995 8732
rect 2995 8676 3051 8732
rect 3051 8676 3055 8732
rect 2991 8672 3055 8676
rect 3071 8732 3135 8736
rect 3071 8676 3075 8732
rect 3075 8676 3131 8732
rect 3131 8676 3135 8732
rect 3071 8672 3135 8676
rect 5269 8732 5333 8736
rect 5269 8676 5273 8732
rect 5273 8676 5329 8732
rect 5329 8676 5333 8732
rect 5269 8672 5333 8676
rect 5349 8732 5413 8736
rect 5349 8676 5353 8732
rect 5353 8676 5409 8732
rect 5409 8676 5413 8732
rect 5349 8672 5413 8676
rect 5429 8732 5493 8736
rect 5429 8676 5433 8732
rect 5433 8676 5489 8732
rect 5489 8676 5493 8732
rect 5429 8672 5493 8676
rect 5509 8732 5573 8736
rect 5509 8676 5513 8732
rect 5513 8676 5569 8732
rect 5569 8676 5573 8732
rect 5509 8672 5573 8676
rect 7707 8732 7771 8736
rect 7707 8676 7711 8732
rect 7711 8676 7767 8732
rect 7767 8676 7771 8732
rect 7707 8672 7771 8676
rect 7787 8732 7851 8736
rect 7787 8676 7791 8732
rect 7791 8676 7847 8732
rect 7847 8676 7851 8732
rect 7787 8672 7851 8676
rect 7867 8732 7931 8736
rect 7867 8676 7871 8732
rect 7871 8676 7927 8732
rect 7927 8676 7931 8732
rect 7867 8672 7931 8676
rect 7947 8732 8011 8736
rect 7947 8676 7951 8732
rect 7951 8676 8007 8732
rect 8007 8676 8011 8732
rect 7947 8672 8011 8676
rect 10145 8732 10209 8736
rect 10145 8676 10149 8732
rect 10149 8676 10205 8732
rect 10205 8676 10209 8732
rect 10145 8672 10209 8676
rect 10225 8732 10289 8736
rect 10225 8676 10229 8732
rect 10229 8676 10285 8732
rect 10285 8676 10289 8732
rect 10225 8672 10289 8676
rect 10305 8732 10369 8736
rect 10305 8676 10309 8732
rect 10309 8676 10365 8732
rect 10365 8676 10369 8732
rect 10305 8672 10369 8676
rect 10385 8732 10449 8736
rect 10385 8676 10389 8732
rect 10389 8676 10445 8732
rect 10445 8676 10449 8732
rect 10385 8672 10449 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 2831 7644 2895 7648
rect 2831 7588 2835 7644
rect 2835 7588 2891 7644
rect 2891 7588 2895 7644
rect 2831 7584 2895 7588
rect 2911 7644 2975 7648
rect 2911 7588 2915 7644
rect 2915 7588 2971 7644
rect 2971 7588 2975 7644
rect 2911 7584 2975 7588
rect 2991 7644 3055 7648
rect 2991 7588 2995 7644
rect 2995 7588 3051 7644
rect 3051 7588 3055 7644
rect 2991 7584 3055 7588
rect 3071 7644 3135 7648
rect 3071 7588 3075 7644
rect 3075 7588 3131 7644
rect 3131 7588 3135 7644
rect 3071 7584 3135 7588
rect 5269 7644 5333 7648
rect 5269 7588 5273 7644
rect 5273 7588 5329 7644
rect 5329 7588 5333 7644
rect 5269 7584 5333 7588
rect 5349 7644 5413 7648
rect 5349 7588 5353 7644
rect 5353 7588 5409 7644
rect 5409 7588 5413 7644
rect 5349 7584 5413 7588
rect 5429 7644 5493 7648
rect 5429 7588 5433 7644
rect 5433 7588 5489 7644
rect 5489 7588 5493 7644
rect 5429 7584 5493 7588
rect 5509 7644 5573 7648
rect 5509 7588 5513 7644
rect 5513 7588 5569 7644
rect 5569 7588 5573 7644
rect 5509 7584 5573 7588
rect 7707 7644 7771 7648
rect 7707 7588 7711 7644
rect 7711 7588 7767 7644
rect 7767 7588 7771 7644
rect 7707 7584 7771 7588
rect 7787 7644 7851 7648
rect 7787 7588 7791 7644
rect 7791 7588 7847 7644
rect 7847 7588 7851 7644
rect 7787 7584 7851 7588
rect 7867 7644 7931 7648
rect 7867 7588 7871 7644
rect 7871 7588 7927 7644
rect 7927 7588 7931 7644
rect 7867 7584 7931 7588
rect 7947 7644 8011 7648
rect 7947 7588 7951 7644
rect 7951 7588 8007 7644
rect 8007 7588 8011 7644
rect 7947 7584 8011 7588
rect 10145 7644 10209 7648
rect 10145 7588 10149 7644
rect 10149 7588 10205 7644
rect 10205 7588 10209 7644
rect 10145 7584 10209 7588
rect 10225 7644 10289 7648
rect 10225 7588 10229 7644
rect 10229 7588 10285 7644
rect 10285 7588 10289 7644
rect 10225 7584 10289 7588
rect 10305 7644 10369 7648
rect 10305 7588 10309 7644
rect 10309 7588 10365 7644
rect 10365 7588 10369 7644
rect 10305 7584 10369 7588
rect 10385 7644 10449 7648
rect 10385 7588 10389 7644
rect 10389 7588 10445 7644
rect 10445 7588 10449 7644
rect 10385 7584 10449 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 2831 6556 2895 6560
rect 2831 6500 2835 6556
rect 2835 6500 2891 6556
rect 2891 6500 2895 6556
rect 2831 6496 2895 6500
rect 2911 6556 2975 6560
rect 2911 6500 2915 6556
rect 2915 6500 2971 6556
rect 2971 6500 2975 6556
rect 2911 6496 2975 6500
rect 2991 6556 3055 6560
rect 2991 6500 2995 6556
rect 2995 6500 3051 6556
rect 3051 6500 3055 6556
rect 2991 6496 3055 6500
rect 3071 6556 3135 6560
rect 3071 6500 3075 6556
rect 3075 6500 3131 6556
rect 3131 6500 3135 6556
rect 3071 6496 3135 6500
rect 5269 6556 5333 6560
rect 5269 6500 5273 6556
rect 5273 6500 5329 6556
rect 5329 6500 5333 6556
rect 5269 6496 5333 6500
rect 5349 6556 5413 6560
rect 5349 6500 5353 6556
rect 5353 6500 5409 6556
rect 5409 6500 5413 6556
rect 5349 6496 5413 6500
rect 5429 6556 5493 6560
rect 5429 6500 5433 6556
rect 5433 6500 5489 6556
rect 5489 6500 5493 6556
rect 5429 6496 5493 6500
rect 5509 6556 5573 6560
rect 5509 6500 5513 6556
rect 5513 6500 5569 6556
rect 5569 6500 5573 6556
rect 5509 6496 5573 6500
rect 7707 6556 7771 6560
rect 7707 6500 7711 6556
rect 7711 6500 7767 6556
rect 7767 6500 7771 6556
rect 7707 6496 7771 6500
rect 7787 6556 7851 6560
rect 7787 6500 7791 6556
rect 7791 6500 7847 6556
rect 7847 6500 7851 6556
rect 7787 6496 7851 6500
rect 7867 6556 7931 6560
rect 7867 6500 7871 6556
rect 7871 6500 7927 6556
rect 7927 6500 7931 6556
rect 7867 6496 7931 6500
rect 7947 6556 8011 6560
rect 7947 6500 7951 6556
rect 7951 6500 8007 6556
rect 8007 6500 8011 6556
rect 7947 6496 8011 6500
rect 10145 6556 10209 6560
rect 10145 6500 10149 6556
rect 10149 6500 10205 6556
rect 10205 6500 10209 6556
rect 10145 6496 10209 6500
rect 10225 6556 10289 6560
rect 10225 6500 10229 6556
rect 10229 6500 10285 6556
rect 10285 6500 10289 6556
rect 10225 6496 10289 6500
rect 10305 6556 10369 6560
rect 10305 6500 10309 6556
rect 10309 6500 10365 6556
rect 10365 6500 10369 6556
rect 10305 6496 10369 6500
rect 10385 6556 10449 6560
rect 10385 6500 10389 6556
rect 10389 6500 10445 6556
rect 10445 6500 10449 6556
rect 10385 6496 10449 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 2831 5468 2895 5472
rect 2831 5412 2835 5468
rect 2835 5412 2891 5468
rect 2891 5412 2895 5468
rect 2831 5408 2895 5412
rect 2911 5468 2975 5472
rect 2911 5412 2915 5468
rect 2915 5412 2971 5468
rect 2971 5412 2975 5468
rect 2911 5408 2975 5412
rect 2991 5468 3055 5472
rect 2991 5412 2995 5468
rect 2995 5412 3051 5468
rect 3051 5412 3055 5468
rect 2991 5408 3055 5412
rect 3071 5468 3135 5472
rect 3071 5412 3075 5468
rect 3075 5412 3131 5468
rect 3131 5412 3135 5468
rect 3071 5408 3135 5412
rect 5269 5468 5333 5472
rect 5269 5412 5273 5468
rect 5273 5412 5329 5468
rect 5329 5412 5333 5468
rect 5269 5408 5333 5412
rect 5349 5468 5413 5472
rect 5349 5412 5353 5468
rect 5353 5412 5409 5468
rect 5409 5412 5413 5468
rect 5349 5408 5413 5412
rect 5429 5468 5493 5472
rect 5429 5412 5433 5468
rect 5433 5412 5489 5468
rect 5489 5412 5493 5468
rect 5429 5408 5493 5412
rect 5509 5468 5573 5472
rect 5509 5412 5513 5468
rect 5513 5412 5569 5468
rect 5569 5412 5573 5468
rect 5509 5408 5573 5412
rect 7707 5468 7771 5472
rect 7707 5412 7711 5468
rect 7711 5412 7767 5468
rect 7767 5412 7771 5468
rect 7707 5408 7771 5412
rect 7787 5468 7851 5472
rect 7787 5412 7791 5468
rect 7791 5412 7847 5468
rect 7847 5412 7851 5468
rect 7787 5408 7851 5412
rect 7867 5468 7931 5472
rect 7867 5412 7871 5468
rect 7871 5412 7927 5468
rect 7927 5412 7931 5468
rect 7867 5408 7931 5412
rect 7947 5468 8011 5472
rect 7947 5412 7951 5468
rect 7951 5412 8007 5468
rect 8007 5412 8011 5468
rect 7947 5408 8011 5412
rect 10145 5468 10209 5472
rect 10145 5412 10149 5468
rect 10149 5412 10205 5468
rect 10205 5412 10209 5468
rect 10145 5408 10209 5412
rect 10225 5468 10289 5472
rect 10225 5412 10229 5468
rect 10229 5412 10285 5468
rect 10285 5412 10289 5468
rect 10225 5408 10289 5412
rect 10305 5468 10369 5472
rect 10305 5412 10309 5468
rect 10309 5412 10365 5468
rect 10365 5412 10369 5468
rect 10305 5408 10369 5412
rect 10385 5468 10449 5472
rect 10385 5412 10389 5468
rect 10389 5412 10445 5468
rect 10445 5412 10449 5468
rect 10385 5408 10449 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 2831 4380 2895 4384
rect 2831 4324 2835 4380
rect 2835 4324 2891 4380
rect 2891 4324 2895 4380
rect 2831 4320 2895 4324
rect 2911 4380 2975 4384
rect 2911 4324 2915 4380
rect 2915 4324 2971 4380
rect 2971 4324 2975 4380
rect 2911 4320 2975 4324
rect 2991 4380 3055 4384
rect 2991 4324 2995 4380
rect 2995 4324 3051 4380
rect 3051 4324 3055 4380
rect 2991 4320 3055 4324
rect 3071 4380 3135 4384
rect 3071 4324 3075 4380
rect 3075 4324 3131 4380
rect 3131 4324 3135 4380
rect 3071 4320 3135 4324
rect 5269 4380 5333 4384
rect 5269 4324 5273 4380
rect 5273 4324 5329 4380
rect 5329 4324 5333 4380
rect 5269 4320 5333 4324
rect 5349 4380 5413 4384
rect 5349 4324 5353 4380
rect 5353 4324 5409 4380
rect 5409 4324 5413 4380
rect 5349 4320 5413 4324
rect 5429 4380 5493 4384
rect 5429 4324 5433 4380
rect 5433 4324 5489 4380
rect 5489 4324 5493 4380
rect 5429 4320 5493 4324
rect 5509 4380 5573 4384
rect 5509 4324 5513 4380
rect 5513 4324 5569 4380
rect 5569 4324 5573 4380
rect 5509 4320 5573 4324
rect 7707 4380 7771 4384
rect 7707 4324 7711 4380
rect 7711 4324 7767 4380
rect 7767 4324 7771 4380
rect 7707 4320 7771 4324
rect 7787 4380 7851 4384
rect 7787 4324 7791 4380
rect 7791 4324 7847 4380
rect 7847 4324 7851 4380
rect 7787 4320 7851 4324
rect 7867 4380 7931 4384
rect 7867 4324 7871 4380
rect 7871 4324 7927 4380
rect 7927 4324 7931 4380
rect 7867 4320 7931 4324
rect 7947 4380 8011 4384
rect 7947 4324 7951 4380
rect 7951 4324 8007 4380
rect 8007 4324 8011 4380
rect 7947 4320 8011 4324
rect 10145 4380 10209 4384
rect 10145 4324 10149 4380
rect 10149 4324 10205 4380
rect 10205 4324 10209 4380
rect 10145 4320 10209 4324
rect 10225 4380 10289 4384
rect 10225 4324 10229 4380
rect 10229 4324 10285 4380
rect 10285 4324 10289 4380
rect 10225 4320 10289 4324
rect 10305 4380 10369 4384
rect 10305 4324 10309 4380
rect 10309 4324 10365 4380
rect 10365 4324 10369 4380
rect 10305 4320 10369 4324
rect 10385 4380 10449 4384
rect 10385 4324 10389 4380
rect 10389 4324 10445 4380
rect 10445 4324 10449 4380
rect 10385 4320 10449 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 2831 3292 2895 3296
rect 2831 3236 2835 3292
rect 2835 3236 2891 3292
rect 2891 3236 2895 3292
rect 2831 3232 2895 3236
rect 2911 3292 2975 3296
rect 2911 3236 2915 3292
rect 2915 3236 2971 3292
rect 2971 3236 2975 3292
rect 2911 3232 2975 3236
rect 2991 3292 3055 3296
rect 2991 3236 2995 3292
rect 2995 3236 3051 3292
rect 3051 3236 3055 3292
rect 2991 3232 3055 3236
rect 3071 3292 3135 3296
rect 3071 3236 3075 3292
rect 3075 3236 3131 3292
rect 3131 3236 3135 3292
rect 3071 3232 3135 3236
rect 5269 3292 5333 3296
rect 5269 3236 5273 3292
rect 5273 3236 5329 3292
rect 5329 3236 5333 3292
rect 5269 3232 5333 3236
rect 5349 3292 5413 3296
rect 5349 3236 5353 3292
rect 5353 3236 5409 3292
rect 5409 3236 5413 3292
rect 5349 3232 5413 3236
rect 5429 3292 5493 3296
rect 5429 3236 5433 3292
rect 5433 3236 5489 3292
rect 5489 3236 5493 3292
rect 5429 3232 5493 3236
rect 5509 3292 5573 3296
rect 5509 3236 5513 3292
rect 5513 3236 5569 3292
rect 5569 3236 5573 3292
rect 5509 3232 5573 3236
rect 7707 3292 7771 3296
rect 7707 3236 7711 3292
rect 7711 3236 7767 3292
rect 7767 3236 7771 3292
rect 7707 3232 7771 3236
rect 7787 3292 7851 3296
rect 7787 3236 7791 3292
rect 7791 3236 7847 3292
rect 7847 3236 7851 3292
rect 7787 3232 7851 3236
rect 7867 3292 7931 3296
rect 7867 3236 7871 3292
rect 7871 3236 7927 3292
rect 7927 3236 7931 3292
rect 7867 3232 7931 3236
rect 7947 3292 8011 3296
rect 7947 3236 7951 3292
rect 7951 3236 8007 3292
rect 8007 3236 8011 3292
rect 7947 3232 8011 3236
rect 10145 3292 10209 3296
rect 10145 3236 10149 3292
rect 10149 3236 10205 3292
rect 10205 3236 10209 3292
rect 10145 3232 10209 3236
rect 10225 3292 10289 3296
rect 10225 3236 10229 3292
rect 10229 3236 10285 3292
rect 10285 3236 10289 3292
rect 10225 3232 10289 3236
rect 10305 3292 10369 3296
rect 10305 3236 10309 3292
rect 10309 3236 10365 3292
rect 10365 3236 10369 3292
rect 10305 3232 10369 3236
rect 10385 3292 10449 3296
rect 10385 3236 10389 3292
rect 10389 3236 10445 3292
rect 10445 3236 10449 3292
rect 10385 3232 10449 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 2831 2204 2895 2208
rect 2831 2148 2835 2204
rect 2835 2148 2891 2204
rect 2891 2148 2895 2204
rect 2831 2144 2895 2148
rect 2911 2204 2975 2208
rect 2911 2148 2915 2204
rect 2915 2148 2971 2204
rect 2971 2148 2975 2204
rect 2911 2144 2975 2148
rect 2991 2204 3055 2208
rect 2991 2148 2995 2204
rect 2995 2148 3051 2204
rect 3051 2148 3055 2204
rect 2991 2144 3055 2148
rect 3071 2204 3135 2208
rect 3071 2148 3075 2204
rect 3075 2148 3131 2204
rect 3131 2148 3135 2204
rect 3071 2144 3135 2148
rect 5269 2204 5333 2208
rect 5269 2148 5273 2204
rect 5273 2148 5329 2204
rect 5329 2148 5333 2204
rect 5269 2144 5333 2148
rect 5349 2204 5413 2208
rect 5349 2148 5353 2204
rect 5353 2148 5409 2204
rect 5409 2148 5413 2204
rect 5349 2144 5413 2148
rect 5429 2204 5493 2208
rect 5429 2148 5433 2204
rect 5433 2148 5489 2204
rect 5489 2148 5493 2204
rect 5429 2144 5493 2148
rect 5509 2204 5573 2208
rect 5509 2148 5513 2204
rect 5513 2148 5569 2204
rect 5569 2148 5573 2204
rect 5509 2144 5573 2148
rect 7707 2204 7771 2208
rect 7707 2148 7711 2204
rect 7711 2148 7767 2204
rect 7767 2148 7771 2204
rect 7707 2144 7771 2148
rect 7787 2204 7851 2208
rect 7787 2148 7791 2204
rect 7791 2148 7847 2204
rect 7847 2148 7851 2204
rect 7787 2144 7851 2148
rect 7867 2204 7931 2208
rect 7867 2148 7871 2204
rect 7871 2148 7927 2204
rect 7927 2148 7931 2204
rect 7867 2144 7931 2148
rect 7947 2204 8011 2208
rect 7947 2148 7951 2204
rect 7951 2148 8007 2204
rect 8007 2148 8011 2204
rect 7947 2144 8011 2148
rect 10145 2204 10209 2208
rect 10145 2148 10149 2204
rect 10149 2148 10205 2204
rect 10205 2148 10209 2204
rect 10145 2144 10209 2148
rect 10225 2204 10289 2208
rect 10225 2148 10229 2204
rect 10229 2148 10285 2204
rect 10285 2148 10289 2204
rect 10225 2144 10289 2148
rect 10305 2204 10369 2208
rect 10305 2148 10309 2204
rect 10309 2148 10365 2204
rect 10365 2148 10369 2204
rect 10305 2144 10369 2148
rect 10385 2204 10449 2208
rect 10385 2148 10389 2204
rect 10389 2148 10445 2204
rect 10445 2148 10449 2204
rect 10385 2144 10449 2148
<< metal4 >>
rect 2163 13632 2483 13648
rect 2163 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2483 13632
rect 2163 12544 2483 13568
rect 2163 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2483 12544
rect 2163 12290 2483 12480
rect 2163 12054 2205 12290
rect 2441 12054 2483 12290
rect 2163 11456 2483 12054
rect 2163 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2483 11456
rect 2163 10368 2483 11392
rect 2163 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2483 10368
rect 2163 9434 2483 10304
rect 2163 9280 2205 9434
rect 2441 9280 2483 9434
rect 2163 9216 2171 9280
rect 2475 9216 2483 9280
rect 2163 9198 2205 9216
rect 2441 9198 2483 9216
rect 2163 8192 2483 9198
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6578 2483 7040
rect 2163 6342 2205 6578
rect 2441 6342 2483 6578
rect 2163 6016 2483 6342
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 3722 2483 3776
rect 2163 3486 2205 3722
rect 2441 3486 2483 3722
rect 2163 2752 2483 3486
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 2823 13088 3143 13648
rect 2823 13024 2831 13088
rect 2895 13024 2911 13088
rect 2975 13024 2991 13088
rect 3055 13024 3071 13088
rect 3135 13024 3143 13088
rect 2823 12950 3143 13024
rect 2823 12714 2865 12950
rect 3101 12714 3143 12950
rect 2823 12000 3143 12714
rect 2823 11936 2831 12000
rect 2895 11936 2911 12000
rect 2975 11936 2991 12000
rect 3055 11936 3071 12000
rect 3135 11936 3143 12000
rect 2823 10912 3143 11936
rect 2823 10848 2831 10912
rect 2895 10848 2911 10912
rect 2975 10848 2991 10912
rect 3055 10848 3071 10912
rect 3135 10848 3143 10912
rect 2823 10094 3143 10848
rect 2823 9858 2865 10094
rect 3101 9858 3143 10094
rect 2823 9824 3143 9858
rect 2823 9760 2831 9824
rect 2895 9760 2911 9824
rect 2975 9760 2991 9824
rect 3055 9760 3071 9824
rect 3135 9760 3143 9824
rect 2823 8736 3143 9760
rect 2823 8672 2831 8736
rect 2895 8672 2911 8736
rect 2975 8672 2991 8736
rect 3055 8672 3071 8736
rect 3135 8672 3143 8736
rect 2823 7648 3143 8672
rect 2823 7584 2831 7648
rect 2895 7584 2911 7648
rect 2975 7584 2991 7648
rect 3055 7584 3071 7648
rect 3135 7584 3143 7648
rect 2823 7238 3143 7584
rect 2823 7002 2865 7238
rect 3101 7002 3143 7238
rect 2823 6560 3143 7002
rect 2823 6496 2831 6560
rect 2895 6496 2911 6560
rect 2975 6496 2991 6560
rect 3055 6496 3071 6560
rect 3135 6496 3143 6560
rect 2823 5472 3143 6496
rect 2823 5408 2831 5472
rect 2895 5408 2911 5472
rect 2975 5408 2991 5472
rect 3055 5408 3071 5472
rect 3135 5408 3143 5472
rect 2823 4384 3143 5408
rect 2823 4320 2831 4384
rect 2895 4382 2911 4384
rect 2975 4382 2991 4384
rect 3055 4382 3071 4384
rect 3135 4320 3143 4384
rect 2823 4146 2865 4320
rect 3101 4146 3143 4320
rect 2823 3296 3143 4146
rect 2823 3232 2831 3296
rect 2895 3232 2911 3296
rect 2975 3232 2991 3296
rect 3055 3232 3071 3296
rect 3135 3232 3143 3296
rect 2823 2208 3143 3232
rect 2823 2144 2831 2208
rect 2895 2144 2911 2208
rect 2975 2144 2991 2208
rect 3055 2144 3071 2208
rect 3135 2144 3143 2208
rect 2823 2128 3143 2144
rect 4601 13632 4921 13648
rect 4601 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4921 13632
rect 4601 12544 4921 13568
rect 4601 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4921 12544
rect 4601 12290 4921 12480
rect 4601 12054 4643 12290
rect 4879 12054 4921 12290
rect 4601 11456 4921 12054
rect 4601 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4921 11456
rect 4601 10368 4921 11392
rect 4601 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4921 10368
rect 4601 9434 4921 10304
rect 4601 9280 4643 9434
rect 4879 9280 4921 9434
rect 4601 9216 4609 9280
rect 4913 9216 4921 9280
rect 4601 9198 4643 9216
rect 4879 9198 4921 9216
rect 4601 8192 4921 9198
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6578 4921 7040
rect 4601 6342 4643 6578
rect 4879 6342 4921 6578
rect 4601 6016 4921 6342
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 3722 4921 3776
rect 4601 3486 4643 3722
rect 4879 3486 4921 3722
rect 4601 2752 4921 3486
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5261 13088 5581 13648
rect 5261 13024 5269 13088
rect 5333 13024 5349 13088
rect 5413 13024 5429 13088
rect 5493 13024 5509 13088
rect 5573 13024 5581 13088
rect 5261 12950 5581 13024
rect 5261 12714 5303 12950
rect 5539 12714 5581 12950
rect 5261 12000 5581 12714
rect 5261 11936 5269 12000
rect 5333 11936 5349 12000
rect 5413 11936 5429 12000
rect 5493 11936 5509 12000
rect 5573 11936 5581 12000
rect 5261 10912 5581 11936
rect 5261 10848 5269 10912
rect 5333 10848 5349 10912
rect 5413 10848 5429 10912
rect 5493 10848 5509 10912
rect 5573 10848 5581 10912
rect 5261 10094 5581 10848
rect 5261 9858 5303 10094
rect 5539 9858 5581 10094
rect 5261 9824 5581 9858
rect 5261 9760 5269 9824
rect 5333 9760 5349 9824
rect 5413 9760 5429 9824
rect 5493 9760 5509 9824
rect 5573 9760 5581 9824
rect 5261 8736 5581 9760
rect 5261 8672 5269 8736
rect 5333 8672 5349 8736
rect 5413 8672 5429 8736
rect 5493 8672 5509 8736
rect 5573 8672 5581 8736
rect 5261 7648 5581 8672
rect 5261 7584 5269 7648
rect 5333 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5581 7648
rect 5261 7238 5581 7584
rect 5261 7002 5303 7238
rect 5539 7002 5581 7238
rect 5261 6560 5581 7002
rect 5261 6496 5269 6560
rect 5333 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5581 6560
rect 5261 5472 5581 6496
rect 5261 5408 5269 5472
rect 5333 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5581 5472
rect 5261 4384 5581 5408
rect 5261 4320 5269 4384
rect 5333 4382 5349 4384
rect 5413 4382 5429 4384
rect 5493 4382 5509 4384
rect 5573 4320 5581 4384
rect 5261 4146 5303 4320
rect 5539 4146 5581 4320
rect 5261 3296 5581 4146
rect 5261 3232 5269 3296
rect 5333 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5581 3296
rect 5261 2208 5581 3232
rect 5261 2144 5269 2208
rect 5333 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5581 2208
rect 5261 2128 5581 2144
rect 7039 13632 7359 13648
rect 7039 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7359 13632
rect 7039 12544 7359 13568
rect 7039 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7359 12544
rect 7039 12290 7359 12480
rect 7039 12054 7081 12290
rect 7317 12054 7359 12290
rect 7039 11456 7359 12054
rect 7039 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7359 11456
rect 7039 10368 7359 11392
rect 7039 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7359 10368
rect 7039 9434 7359 10304
rect 7039 9280 7081 9434
rect 7317 9280 7359 9434
rect 7039 9216 7047 9280
rect 7351 9216 7359 9280
rect 7039 9198 7081 9216
rect 7317 9198 7359 9216
rect 7039 8192 7359 9198
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6578 7359 7040
rect 7039 6342 7081 6578
rect 7317 6342 7359 6578
rect 7039 6016 7359 6342
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 3722 7359 3776
rect 7039 3486 7081 3722
rect 7317 3486 7359 3722
rect 7039 2752 7359 3486
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 7699 13088 8019 13648
rect 7699 13024 7707 13088
rect 7771 13024 7787 13088
rect 7851 13024 7867 13088
rect 7931 13024 7947 13088
rect 8011 13024 8019 13088
rect 7699 12950 8019 13024
rect 7699 12714 7741 12950
rect 7977 12714 8019 12950
rect 7699 12000 8019 12714
rect 7699 11936 7707 12000
rect 7771 11936 7787 12000
rect 7851 11936 7867 12000
rect 7931 11936 7947 12000
rect 8011 11936 8019 12000
rect 7699 10912 8019 11936
rect 7699 10848 7707 10912
rect 7771 10848 7787 10912
rect 7851 10848 7867 10912
rect 7931 10848 7947 10912
rect 8011 10848 8019 10912
rect 7699 10094 8019 10848
rect 7699 9858 7741 10094
rect 7977 9858 8019 10094
rect 7699 9824 8019 9858
rect 7699 9760 7707 9824
rect 7771 9760 7787 9824
rect 7851 9760 7867 9824
rect 7931 9760 7947 9824
rect 8011 9760 8019 9824
rect 7699 8736 8019 9760
rect 7699 8672 7707 8736
rect 7771 8672 7787 8736
rect 7851 8672 7867 8736
rect 7931 8672 7947 8736
rect 8011 8672 8019 8736
rect 7699 7648 8019 8672
rect 7699 7584 7707 7648
rect 7771 7584 7787 7648
rect 7851 7584 7867 7648
rect 7931 7584 7947 7648
rect 8011 7584 8019 7648
rect 7699 7238 8019 7584
rect 7699 7002 7741 7238
rect 7977 7002 8019 7238
rect 7699 6560 8019 7002
rect 7699 6496 7707 6560
rect 7771 6496 7787 6560
rect 7851 6496 7867 6560
rect 7931 6496 7947 6560
rect 8011 6496 8019 6560
rect 7699 5472 8019 6496
rect 7699 5408 7707 5472
rect 7771 5408 7787 5472
rect 7851 5408 7867 5472
rect 7931 5408 7947 5472
rect 8011 5408 8019 5472
rect 7699 4384 8019 5408
rect 7699 4320 7707 4384
rect 7771 4382 7787 4384
rect 7851 4382 7867 4384
rect 7931 4382 7947 4384
rect 8011 4320 8019 4384
rect 7699 4146 7741 4320
rect 7977 4146 8019 4320
rect 7699 3296 8019 4146
rect 7699 3232 7707 3296
rect 7771 3232 7787 3296
rect 7851 3232 7867 3296
rect 7931 3232 7947 3296
rect 8011 3232 8019 3296
rect 7699 2208 8019 3232
rect 7699 2144 7707 2208
rect 7771 2144 7787 2208
rect 7851 2144 7867 2208
rect 7931 2144 7947 2208
rect 8011 2144 8019 2208
rect 7699 2128 8019 2144
rect 9477 13632 9797 13648
rect 9477 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9797 13632
rect 9477 12544 9797 13568
rect 9477 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9797 12544
rect 9477 12290 9797 12480
rect 9477 12054 9519 12290
rect 9755 12054 9797 12290
rect 9477 11456 9797 12054
rect 9477 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9797 11456
rect 9477 10368 9797 11392
rect 9477 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9797 10368
rect 9477 9434 9797 10304
rect 9477 9280 9519 9434
rect 9755 9280 9797 9434
rect 9477 9216 9485 9280
rect 9789 9216 9797 9280
rect 9477 9198 9519 9216
rect 9755 9198 9797 9216
rect 9477 8192 9797 9198
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6578 9797 7040
rect 9477 6342 9519 6578
rect 9755 6342 9797 6578
rect 9477 6016 9797 6342
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 3722 9797 3776
rect 9477 3486 9519 3722
rect 9755 3486 9797 3722
rect 9477 2752 9797 3486
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10137 13088 10457 13648
rect 10137 13024 10145 13088
rect 10209 13024 10225 13088
rect 10289 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10457 13088
rect 10137 12950 10457 13024
rect 10137 12714 10179 12950
rect 10415 12714 10457 12950
rect 10137 12000 10457 12714
rect 10137 11936 10145 12000
rect 10209 11936 10225 12000
rect 10289 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10457 12000
rect 10137 10912 10457 11936
rect 10137 10848 10145 10912
rect 10209 10848 10225 10912
rect 10289 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10457 10912
rect 10137 10094 10457 10848
rect 10137 9858 10179 10094
rect 10415 9858 10457 10094
rect 10137 9824 10457 9858
rect 10137 9760 10145 9824
rect 10209 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10457 9824
rect 10137 8736 10457 9760
rect 10137 8672 10145 8736
rect 10209 8672 10225 8736
rect 10289 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10457 8736
rect 10137 7648 10457 8672
rect 10137 7584 10145 7648
rect 10209 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10457 7648
rect 10137 7238 10457 7584
rect 10137 7002 10179 7238
rect 10415 7002 10457 7238
rect 10137 6560 10457 7002
rect 10137 6496 10145 6560
rect 10209 6496 10225 6560
rect 10289 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10457 6560
rect 10137 5472 10457 6496
rect 10137 5408 10145 5472
rect 10209 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10457 5472
rect 10137 4384 10457 5408
rect 10137 4320 10145 4384
rect 10209 4382 10225 4384
rect 10289 4382 10305 4384
rect 10369 4382 10385 4384
rect 10449 4320 10457 4384
rect 10137 4146 10179 4320
rect 10415 4146 10457 4320
rect 10137 3296 10457 4146
rect 10137 3232 10145 3296
rect 10209 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10457 3296
rect 10137 2208 10457 3232
rect 10137 2144 10145 2208
rect 10209 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10457 2208
rect 10137 2128 10457 2144
<< via4 >>
rect 2205 12054 2441 12290
rect 2205 9280 2441 9434
rect 2205 9216 2235 9280
rect 2235 9216 2251 9280
rect 2251 9216 2315 9280
rect 2315 9216 2331 9280
rect 2331 9216 2395 9280
rect 2395 9216 2411 9280
rect 2411 9216 2441 9280
rect 2205 9198 2441 9216
rect 2205 6342 2441 6578
rect 2205 3486 2441 3722
rect 2865 12714 3101 12950
rect 2865 9858 3101 10094
rect 2865 7002 3101 7238
rect 2865 4320 2895 4382
rect 2895 4320 2911 4382
rect 2911 4320 2975 4382
rect 2975 4320 2991 4382
rect 2991 4320 3055 4382
rect 3055 4320 3071 4382
rect 3071 4320 3101 4382
rect 2865 4146 3101 4320
rect 4643 12054 4879 12290
rect 4643 9280 4879 9434
rect 4643 9216 4673 9280
rect 4673 9216 4689 9280
rect 4689 9216 4753 9280
rect 4753 9216 4769 9280
rect 4769 9216 4833 9280
rect 4833 9216 4849 9280
rect 4849 9216 4879 9280
rect 4643 9198 4879 9216
rect 4643 6342 4879 6578
rect 4643 3486 4879 3722
rect 5303 12714 5539 12950
rect 5303 9858 5539 10094
rect 5303 7002 5539 7238
rect 5303 4320 5333 4382
rect 5333 4320 5349 4382
rect 5349 4320 5413 4382
rect 5413 4320 5429 4382
rect 5429 4320 5493 4382
rect 5493 4320 5509 4382
rect 5509 4320 5539 4382
rect 5303 4146 5539 4320
rect 7081 12054 7317 12290
rect 7081 9280 7317 9434
rect 7081 9216 7111 9280
rect 7111 9216 7127 9280
rect 7127 9216 7191 9280
rect 7191 9216 7207 9280
rect 7207 9216 7271 9280
rect 7271 9216 7287 9280
rect 7287 9216 7317 9280
rect 7081 9198 7317 9216
rect 7081 6342 7317 6578
rect 7081 3486 7317 3722
rect 7741 12714 7977 12950
rect 7741 9858 7977 10094
rect 7741 7002 7977 7238
rect 7741 4320 7771 4382
rect 7771 4320 7787 4382
rect 7787 4320 7851 4382
rect 7851 4320 7867 4382
rect 7867 4320 7931 4382
rect 7931 4320 7947 4382
rect 7947 4320 7977 4382
rect 7741 4146 7977 4320
rect 9519 12054 9755 12290
rect 9519 9280 9755 9434
rect 9519 9216 9549 9280
rect 9549 9216 9565 9280
rect 9565 9216 9629 9280
rect 9629 9216 9645 9280
rect 9645 9216 9709 9280
rect 9709 9216 9725 9280
rect 9725 9216 9755 9280
rect 9519 9198 9755 9216
rect 9519 6342 9755 6578
rect 9519 3486 9755 3722
rect 10179 12714 10415 12950
rect 10179 9858 10415 10094
rect 10179 7002 10415 7238
rect 10179 4320 10209 4382
rect 10209 4320 10225 4382
rect 10225 4320 10289 4382
rect 10289 4320 10305 4382
rect 10305 4320 10369 4382
rect 10369 4320 10385 4382
rect 10385 4320 10415 4382
rect 10179 4146 10415 4320
<< metal5 >>
rect 1056 12950 10904 12992
rect 1056 12714 2865 12950
rect 3101 12714 5303 12950
rect 5539 12714 7741 12950
rect 7977 12714 10179 12950
rect 10415 12714 10904 12950
rect 1056 12672 10904 12714
rect 1056 12290 10904 12332
rect 1056 12054 2205 12290
rect 2441 12054 4643 12290
rect 4879 12054 7081 12290
rect 7317 12054 9519 12290
rect 9755 12054 10904 12290
rect 1056 12012 10904 12054
rect 1056 10094 10904 10136
rect 1056 9858 2865 10094
rect 3101 9858 5303 10094
rect 5539 9858 7741 10094
rect 7977 9858 10179 10094
rect 10415 9858 10904 10094
rect 1056 9816 10904 9858
rect 1056 9434 10904 9476
rect 1056 9198 2205 9434
rect 2441 9198 4643 9434
rect 4879 9198 7081 9434
rect 7317 9198 9519 9434
rect 9755 9198 10904 9434
rect 1056 9156 10904 9198
rect 1056 7238 10904 7280
rect 1056 7002 2865 7238
rect 3101 7002 5303 7238
rect 5539 7002 7741 7238
rect 7977 7002 10179 7238
rect 10415 7002 10904 7238
rect 1056 6960 10904 7002
rect 1056 6578 10904 6620
rect 1056 6342 2205 6578
rect 2441 6342 4643 6578
rect 4879 6342 7081 6578
rect 7317 6342 9519 6578
rect 9755 6342 10904 6578
rect 1056 6300 10904 6342
rect 1056 4382 10904 4424
rect 1056 4146 2865 4382
rect 3101 4146 5303 4382
rect 5539 4146 7741 4382
rect 7977 4146 10179 4382
rect 10415 4146 10904 4382
rect 1056 4104 10904 4146
rect 1056 3722 10904 3764
rect 1056 3486 2205 3722
rect 2441 3486 4643 3722
rect 4879 3486 7081 3722
rect 7317 3486 9519 3722
rect 9755 3486 10904 3722
rect 1056 3444 10904 3486
use sky130_fd_sc_hd__or2_1  _161_
timestamp 0
transform 1 0 1748 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _162_
timestamp 0
transform 1 0 2208 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _163_
timestamp 0
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 0
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _165_
timestamp 0
transform 1 0 3036 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _166_
timestamp 0
transform 1 0 3128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _167_
timestamp 0
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _168_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _169_
timestamp 0
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _170_
timestamp 0
transform 1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _171_
timestamp 0
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _172_
timestamp 0
transform 1 0 6808 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _173_
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _174_
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _175_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _176_
timestamp 0
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _177_
timestamp 0
transform 1 0 5888 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _178_
timestamp 0
transform -1 0 7176 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _179_
timestamp 0
transform -1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _180_
timestamp 0
transform 1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _181_
timestamp 0
transform -1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _182_
timestamp 0
transform 1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _183_
timestamp 0
transform 1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _184_
timestamp 0
transform -1 0 7544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 0
transform -1 0 8004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _186_
timestamp 0
transform -1 0 4508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _187_
timestamp 0
transform 1 0 6256 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _188_
timestamp 0
transform -1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _189_
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _190_
timestamp 0
transform -1 0 8280 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _191_
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _192_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _193_
timestamp 0
transform 1 0 9200 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _194_
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _195_
timestamp 0
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _196_
timestamp 0
transform 1 0 7912 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _197_
timestamp 0
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _198_
timestamp 0
transform 1 0 8648 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _199_
timestamp 0
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _200_
timestamp 0
transform 1 0 9108 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 0
transform -1 0 10212 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 0
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _203_
timestamp 0
transform 1 0 9476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_
timestamp 0
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 0
transform -1 0 8648 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _206_
timestamp 0
transform -1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _207_
timestamp 0
transform 1 0 7544 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _208_
timestamp 0
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _209_
timestamp 0
transform 1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _210_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _211_
timestamp 0
transform -1 0 9660 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 0
transform 1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _213_
timestamp 0
transform -1 0 2760 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _214_
timestamp 0
transform 1 0 1564 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _215_
timestamp 0
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _216_
timestamp 0
transform 1 0 1656 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _217_
timestamp 0
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _218_
timestamp 0
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _219_
timestamp 0
transform 1 0 2668 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _220_
timestamp 0
transform 1 0 1932 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _221_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _222_
timestamp 0
transform -1 0 3036 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__o41a_1  _223_
timestamp 0
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _225_
timestamp 0
transform 1 0 1840 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _227_
timestamp 0
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _228_
timestamp 0
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _229_
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _230_
timestamp 0
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _231_
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _232_
timestamp 0
transform 1 0 2392 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _233_
timestamp 0
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _234_
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 0
transform -1 0 3404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _236_
timestamp 0
transform -1 0 3864 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 0
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _238_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _239_
timestamp 0
transform -1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _240_
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _241_
timestamp 0
transform 1 0 3864 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _242_
timestamp 0
transform 1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _243_
timestamp 0
transform 1 0 1748 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _244_
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _245_
timestamp 0
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _246_
timestamp 0
transform 1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _247_
timestamp 0
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_2  _248_
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _249_
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 0
transform 1 0 2208 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 0
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _252_
timestamp 0
transform -1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _253_
timestamp 0
transform 1 0 4876 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_1  _254_
timestamp 0
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _255_
timestamp 0
transform -1 0 2484 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _256_
timestamp 0
transform 1 0 2024 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _257_
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 0
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_2  _260_
timestamp 0
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _261_
timestamp 0
transform -1 0 4968 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _262_
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _263_
timestamp 0
transform -1 0 5520 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _264_
timestamp 0
transform 1 0 6440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _265_
timestamp 0
transform 1 0 7360 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _266_
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _267_
timestamp 0
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _268_
timestamp 0
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _269_
timestamp 0
transform 1 0 7912 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _270_
timestamp 0
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _271_
timestamp 0
transform 1 0 2852 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _272_
timestamp 0
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _273_
timestamp 0
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _274_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp 0
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 0
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _277_
timestamp 0
transform -1 0 6624 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 0
transform -1 0 2944 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _279_
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _280_
timestamp 0
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _281_
timestamp 0
transform 1 0 5152 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _282_
timestamp 0
transform 1 0 5520 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _283_
timestamp 0
transform 1 0 7544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _284_
timestamp 0
transform -1 0 7084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _285_
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 0
transform -1 0 7268 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _287_
timestamp 0
transform -1 0 7912 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 0
transform -1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _289_
timestamp 0
transform 1 0 6440 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _290_
timestamp 0
transform -1 0 5244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _291_
timestamp 0
transform -1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _292_
timestamp 0
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 0
transform -1 0 5796 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _294_
timestamp 0
transform 1 0 6992 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _295_
timestamp 0
transform 1 0 6532 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _296_
timestamp 0
transform -1 0 8556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _297_
timestamp 0
transform -1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _298_
timestamp 0
transform 1 0 6808 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _299_
timestamp 0
transform -1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _300_
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _301_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _302_
timestamp 0
transform 1 0 6072 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _303_
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _304_
timestamp 0
transform -1 0 10304 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _305_
timestamp 0
transform 1 0 4232 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _306_
timestamp 0
transform -1 0 5704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _307_
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _308_
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _309_
timestamp 0
transform -1 0 5152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _310_
timestamp 0
transform -1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _311_
timestamp 0
transform -1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _312_
timestamp 0
transform 1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 0
transform -1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _314_
timestamp 0
transform -1 0 5244 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _315_
timestamp 0
transform -1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _316_
timestamp 0
transform 1 0 5704 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _317_
timestamp 0
transform -1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _318_
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _319_
timestamp 0
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _320_
timestamp 0
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _321_
timestamp 0
transform 1 0 9476 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _322_
timestamp 0
transform 1 0 3956 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _323_
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _324_
timestamp 0
transform -1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _325_
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _326_
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _327_
timestamp 0
transform -1 0 4692 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _328_
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 0
transform -1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_10
timestamp 0
transform 1 0 2024 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_18
timestamp 0
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_31
timestamp 0
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_42
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49
timestamp 0
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_71
timestamp 0
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_75
timestamp 0
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_80
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_92
timestamp 0
transform 1 0 9568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_100
timestamp 0
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_7
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_17
timestamp 0
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 0
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_38
timestamp 0
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 0
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_91
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_6
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_26
timestamp 0
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_31
timestamp 0
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_65
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_91
timestamp 0
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 0
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_18
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_24
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_34
timestamp 0
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 0
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_60
timestamp 0
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_72
timestamp 0
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_24
timestamp 0
transform 1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_73
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_85
timestamp 0
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_49
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_66
timestamp 0
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_31
timestamp 0
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_61
timestamp 0
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_98
timestamp 0
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_102
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_57
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_70
timestamp 0
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 0
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_88
timestamp 0
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_99
timestamp 0
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_20
timestamp 0
transform 1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_28
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_46
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_51
timestamp 0
transform 1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_59
timestamp 0
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_76
timestamp 0
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_13
timestamp 0
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_25
timestamp 0
transform 1 0 3404 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_33
timestamp 0
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_52
timestamp 0
transform 1 0 5888 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_82
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_97
timestamp 0
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 0
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_45
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 0
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_34
timestamp 0
transform 1 0 4232 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_46
timestamp 0
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_64
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_76
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_80
timestamp 0
transform 1 0 8464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_98
timestamp 0
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_102
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_11
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 0
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_37
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_43
timestamp 0
transform 1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_50
timestamp 0
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_62
timestamp 0
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_91
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_9
timestamp 0
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 0
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_33
timestamp 0
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_78
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_90
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_98
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_6
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_17
timestamp 0
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_49
timestamp 0
transform 1 0 5612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_55
timestamp 0
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_61
timestamp 0
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_70
timestamp 0
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_100
timestamp 0
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_17
timestamp 0
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_44
timestamp 0
transform 1 0 5152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 0
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_95
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 0
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_25
timestamp 0
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_37
timestamp 0
transform 1 0 4508 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_67
timestamp 0
transform 1 0 7268 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_79
timestamp 0
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_91
timestamp 0
transform 1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 0
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 0
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 0
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 0
transform 1 0 3036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 0
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 0
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 0
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 0
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 0
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 0
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_21
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_22
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_23
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_24
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_25
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_26
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_27
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_28
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_29
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_30
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_31
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_32
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_33
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_34
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_35
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_36
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_37
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_38
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_39
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_40
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_41
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_44
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_49
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_50
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_51
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_52
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_53
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_54
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_55
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_56
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_57
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_58
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_59
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_60
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_61
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_62
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_63
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_64
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_65
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_66
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_67
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_68
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_69
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_70
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_71
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_72
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_73
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_74
timestamp 0
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_75
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5980 13056 5980 13056 4 VGND
rlabel metal1 s 5980 13600 5980 13600 4 VPWR
rlabel metal3 s 0 6264 800 6384 4 A[0]
port 1 nsew
rlabel metal3 s 1050 5508 1050 5508 4 A[1]
rlabel metal3 s 0 4632 800 4752 4 A[2]
port 3 nsew
rlabel metal3 s 0 3816 800 3936 4 A[3]
port 4 nsew
rlabel metal3 s 0 3000 800 3120 4 A[4]
port 5 nsew
rlabel metal3 s 0 2184 800 2304 4 A[5]
port 6 nsew
rlabel metal3 s 1096 1428 1096 1428 4 A[6]
rlabel metal3 s 1234 612 1234 612 4 A[7]
rlabel metal3 s 1694 12852 1694 12852 4 B[0]
rlabel metal3 s 1188 12036 1188 12036 4 B[1]
rlabel metal3 s 0 11160 800 11280 4 B[2]
port 11 nsew
rlabel metal3 s 0 10344 800 10464 4 B[3]
port 12 nsew
rlabel metal3 s 1096 9588 1096 9588 4 B[4]
rlabel metal3 s 0 8712 800 8832 4 B[5]
port 14 nsew
rlabel metal3 s 1050 7956 1050 7956 4 B[6]
rlabel metal3 s 0 7080 800 7200 4 B[7]
port 16 nsew
rlabel metal2 s 4370 8364 4370 8364 4 _000_
rlabel metal1 s 3588 11866 3588 11866 4 _001_
rlabel metal2 s 3450 11424 3450 11424 4 _002_
rlabel metal1 s 4554 11730 4554 11730 4 _003_
rlabel metal1 s 5198 12954 5198 12954 4 _004_
rlabel metal2 s 4186 11900 4186 11900 4 _005_
rlabel metal1 s 4968 11594 4968 11594 4 _006_
rlabel metal1 s 4278 10574 4278 10574 4 _007_
rlabel metal1 s 4738 11084 4738 11084 4 _008_
rlabel metal2 s 2070 9724 2070 9724 4 _009_
rlabel metal1 s 3772 8466 3772 8466 4 _010_
rlabel metal2 s 4186 7616 4186 7616 4 _011_
rlabel metal1 s 4830 8296 4830 8296 4 _012_
rlabel metal1 s 4186 6426 4186 6426 4 _013_
rlabel metal2 s 4922 7276 4922 7276 4 _014_
rlabel metal2 s 4278 6970 4278 6970 4 _015_
rlabel metal1 s 5014 5100 5014 5100 4 _016_
rlabel metal1 s 2622 11016 2622 11016 4 _017_
rlabel metal1 s 5106 11322 5106 11322 4 _018_
rlabel metal1 s 4922 5168 4922 5168 4 _019_
rlabel metal1 s 5658 5304 5658 5304 4 _020_
rlabel metal1 s 2300 7174 2300 7174 4 _021_
rlabel metal2 s 2622 3162 2622 3162 4 _022_
rlabel metal2 s 3634 3196 3634 3196 4 _023_
rlabel metal1 s 4830 4080 4830 4080 4 _024_
rlabel metal1 s 4922 4658 4922 4658 4 _025_
rlabel metal1 s 4968 3638 4968 3638 4 _026_
rlabel metal1 s 5106 4114 5106 4114 4 _027_
rlabel metal2 s 5474 3706 5474 3706 4 _028_
rlabel metal1 s 8832 3502 8832 3502 4 _029_
rlabel metal1 s 7406 5678 7406 5678 4 _030_
rlabel metal2 s 7590 4879 7590 4879 4 _031_
rlabel metal2 s 8142 5151 8142 5151 4 _032_
rlabel metal2 s 8142 3706 8142 3706 4 _033_
rlabel metal1 s 7866 4080 7866 4080 4 _034_
rlabel metal2 s 8418 3196 8418 3196 4 _035_
rlabel metal1 s 3174 4046 3174 4046 4 _036_
rlabel metal1 s 2714 4080 2714 4080 4 _037_
rlabel metal2 s 3266 3638 3266 3638 4 _038_
rlabel metal1 s 8605 3162 8605 3162 4 _039_
rlabel metal1 s 4094 2992 4094 2992 4 _040_
rlabel metal2 s 4738 3332 4738 3332 4 _041_
rlabel metal2 s 6026 3264 6026 3264 4 _042_
rlabel metal1 s 4738 2958 4738 2958 4 _043_
rlabel metal2 s 5198 3298 5198 3298 4 _044_
rlabel metal1 s 5336 3706 5336 3706 4 _045_
rlabel metal1 s 5658 3162 5658 3162 4 _046_
rlabel metal1 s 6762 3060 6762 3060 4 _047_
rlabel metal2 s 7682 3706 7682 3706 4 _048_
rlabel metal2 s 7406 3706 7406 3706 4 _049_
rlabel metal1 s 6992 3162 6992 3162 4 _050_
rlabel metal1 s 7314 3536 7314 3536 4 _051_
rlabel metal2 s 6854 3196 6854 3196 4 _052_
rlabel metal1 s 6946 3060 6946 3060 4 _053_
rlabel metal2 s 5106 12002 5106 12002 4 _054_
rlabel metal2 s 5658 11900 5658 11900 4 _055_
rlabel metal1 s 5382 12750 5382 12750 4 _056_
rlabel metal1 s 7268 12614 7268 12614 4 _057_
rlabel metal2 s 6578 12036 6578 12036 4 _058_
rlabel metal1 s 8878 12070 8878 12070 4 _059_
rlabel metal1 s 7038 12172 7038 12172 4 _060_
rlabel metal1 s 6808 12614 6808 12614 4 _061_
rlabel metal1 s 5198 11152 5198 11152 4 _062_
rlabel metal1 s 5980 11322 5980 11322 4 _063_
rlabel metal1 s 6808 12342 6808 12342 4 _064_
rlabel metal2 s 9890 11288 9890 11288 4 _065_
rlabel metal1 s 8972 11186 8972 11186 4 _066_
rlabel metal1 s 4784 10506 4784 10506 4 _067_
rlabel metal2 s 5842 10438 5842 10438 4 _068_
rlabel metal1 s 5382 10608 5382 10608 4 _069_
rlabel metal1 s 4738 10778 4738 10778 4 _070_
rlabel metal1 s 6072 11254 6072 11254 4 _071_
rlabel metal1 s 9844 8466 9844 8466 4 _072_
rlabel metal2 s 5014 8092 5014 8092 4 _073_
rlabel metal1 s 5658 7242 5658 7242 4 _074_
rlabel metal1 s 5474 7820 5474 7820 4 _075_
rlabel metal1 s 6072 6154 6072 6154 4 _076_
rlabel metal1 s 5106 6800 5106 6800 4 _077_
rlabel metal1 s 5704 6970 5704 6970 4 _078_
rlabel metal1 s 5566 8058 5566 8058 4 _079_
rlabel metal1 s 9292 8466 9292 8466 4 _080_
rlabel metal2 s 10074 6494 10074 6494 4 _081_
rlabel metal2 s 3910 7548 3910 7548 4 _082_
rlabel metal2 s 4462 7038 4462 7038 4 _083_
rlabel metal1 s 1978 6868 1978 6868 4 _084_
rlabel metal1 s 2622 6732 2622 6732 4 _085_
rlabel metal1 s 4186 6698 4186 6698 4 _086_
rlabel metal1 s 8602 6698 8602 6698 4 _087_
rlabel metal1 s 9844 6766 9844 6766 4 _088_
rlabel metal1 s 2400 11050 2400 11050 4 _089_
rlabel metal2 s 2530 4726 2530 4726 4 _090_
rlabel metal2 s 9016 8466 9016 8466 4 _091_
rlabel metal2 s 1978 11832 1978 11832 4 _092_
rlabel metal1 s 9844 11322 9844 11322 4 _093_
rlabel metal1 s 10028 9554 10028 9554 4 _094_
rlabel metal1 s 7590 6324 7590 6324 4 _095_
rlabel metal2 s 6946 9214 6946 9214 4 _096_
rlabel metal1 s 3220 9078 3220 9078 4 _097_
rlabel metal1 s 6670 8874 6670 8874 4 _098_
rlabel metal1 s 2622 9520 2622 9520 4 _099_
rlabel metal1 s 7774 7888 7774 7888 4 _100_
rlabel metal1 s 7682 11322 7682 11322 4 _101_
rlabel metal1 s 7528 8534 7528 8534 4 _102_
rlabel metal1 s 8740 8262 8740 8262 4 _103_
rlabel metal1 s 6302 8534 6302 8534 4 _104_
rlabel metal2 s 6946 8109 6946 8109 4 _105_
rlabel metal1 s 7498 7820 7498 7820 4 _106_
rlabel metal1 s 7774 6766 7774 6766 4 _107_
rlabel metal2 s 7498 7242 7498 7242 4 _108_
rlabel metal2 s 7498 6426 7498 6426 4 _109_
rlabel metal1 s 9062 6222 9062 6222 4 _110_
rlabel metal1 s 9752 9486 9752 9486 4 _111_
rlabel metal1 s 7544 8602 7544 8602 4 _112_
rlabel metal2 s 8786 9350 8786 9350 4 _113_
rlabel metal2 s 3910 10914 3910 10914 4 _114_
rlabel metal1 s 7590 12818 7590 12818 4 _115_
rlabel metal1 s 8096 11254 8096 11254 4 _116_
rlabel metal1 s 7958 11016 7958 11016 4 _117_
rlabel metal2 s 8970 10268 8970 10268 4 _118_
rlabel metal1 s 9154 9452 9154 9452 4 _119_
rlabel metal2 s 9706 9724 9706 9724 4 _120_
rlabel metal1 s 9200 6766 9200 6766 4 _121_
rlabel metal1 s 9798 6290 9798 6290 4 _122_
rlabel metal1 s 8234 11764 8234 11764 4 _123_
rlabel metal2 s 8418 11492 8418 11492 4 _124_
rlabel metal1 s 9062 11696 9062 11696 4 _125_
rlabel metal2 s 10258 11526 10258 11526 4 _126_
rlabel metal2 s 9338 9146 9338 9146 4 _127_
rlabel metal1 s 9844 8942 9844 8942 4 _128_
rlabel metal1 s 10028 8466 10028 8466 4 _129_
rlabel metal2 s 8694 6154 8694 6154 4 _130_
rlabel metal1 s 9476 5202 9476 5202 4 _131_
rlabel metal2 s 8418 6596 8418 6596 4 _132_
rlabel metal1 s 8004 8466 8004 8466 4 _133_
rlabel metal1 s 7958 8398 7958 8398 4 _134_
rlabel metal1 s 8188 6834 8188 6834 4 _135_
rlabel metal2 s 8510 5882 8510 5882 4 _136_
rlabel metal1 s 8924 5678 8924 5678 4 _137_
rlabel metal2 s 9338 5338 9338 5338 4 _138_
rlabel metal1 s 7866 5202 7866 5202 4 _139_
rlabel metal2 s 2438 12835 2438 12835 4 _140_
rlabel metal2 s 5474 6817 5474 6817 4 _141_
rlabel metal1 s 2668 12750 2668 12750 4 _142_
rlabel metal2 s 2990 6817 2990 6817 4 _143_
rlabel metal2 s 2254 13124 2254 13124 4 _144_
rlabel metal1 s 1978 13158 1978 13158 4 _145_
rlabel metal1 s 1886 5100 1886 5100 4 _146_
rlabel metal1 s 2668 5202 2668 5202 4 _147_
rlabel metal1 s 4278 5202 4278 5202 4 _148_
rlabel metal1 s 5842 5168 5842 5168 4 _149_
rlabel metal2 s 2714 12036 2714 12036 4 _150_
rlabel metal2 s 2070 8398 2070 8398 4 _151_
rlabel metal1 s 2346 5746 2346 5746 4 _152_
rlabel metal2 s 3818 5032 3818 5032 4 _153_
rlabel metal1 s 4738 4522 4738 4522 4 _154_
rlabel metal1 s 3634 4250 3634 4250 4 _155_
rlabel metal2 s 4370 4998 4370 4998 4 _156_
rlabel metal1 s 2622 7344 2622 7344 4 _157_
rlabel metal1 s 4370 6358 4370 6358 4 _158_
rlabel metal1 s 2070 9418 2070 9418 4 _159_
rlabel metal2 s 3910 9316 3910 9316 4 _160_
rlabel metal2 s 1610 6528 1610 6528 4 net1
rlabel metal1 s 6532 11118 6532 11118 4 net10
rlabel metal1 s 2530 11152 2530 11152 4 net11
rlabel metal2 s 1978 10030 1978 10030 4 net12
rlabel metal1 s 2162 8024 2162 8024 4 net13
rlabel metal1 s 2392 7854 2392 7854 4 net14
rlabel metal1 s 2346 7310 2346 7310 4 net15
rlabel metal1 s 2622 7208 2622 7208 4 net16
rlabel metal2 s 3358 12988 3358 12988 4 net17
rlabel metal2 s 2806 12716 2806 12716 4 net18
rlabel metal1 s 2714 12852 2714 12852 4 net19
rlabel metal2 s 7314 6222 7314 6222 4 net2
rlabel metal2 s 8602 12988 8602 12988 4 net20
rlabel metal3 s 6118 12325 6118 12325 4 net21
rlabel metal1 s 10166 10642 10166 10642 4 net22
rlabel metal1 s 10258 8432 10258 8432 4 net23
rlabel metal2 s 10258 7174 10258 7174 4 net24
rlabel metal1 s 7958 4998 7958 4998 4 net25
rlabel metal1 s 10258 3570 10258 3570 4 net26
rlabel metal1 s 8832 2822 8832 2822 4 net27
rlabel metal1 s 4554 8908 4554 8908 4 net3
rlabel metal2 s 1610 3774 1610 3774 4 net4
rlabel metal1 s 1748 6766 1748 6766 4 net5
rlabel metal1 s 2024 5270 2024 5270 4 net6
rlabel metal2 s 3910 3247 3910 3247 4 net7
rlabel metal2 s 6394 3281 6394 3281 4 net8
rlabel metal1 s 3266 13226 3266 13226 4 net9
rlabel metal3 s 2154 15300 2154 15300 4 opcode[0]
rlabel metal3 s 1050 14484 1050 14484 4 opcode[1]
rlabel metal3 s 1119 13668 1119 13668 4 opcode[2]
rlabel metal2 s 10442 13991 10442 13991 4 out[0]
rlabel metal3 s 10442 12597 10442 12597 4 out[1]
rlabel metal2 s 10442 10727 10442 10727 4 out[2]
rlabel metal1 s 10672 8602 10672 8602 4 out[3]
rlabel metal2 s 10442 7021 10442 7021 4 out[4]
rlabel metal3 s 10442 4981 10442 4981 4 out[5]
rlabel metal1 s 10488 3366 10488 3366 4 out[6]
rlabel metal1 s 10028 2278 10028 2278 4 out[7]
flabel metal3 s 400 6324 400 6324 0 FreeSans 600 0 0 0 A[0]
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 A[1]
port 2 nsew
flabel metal3 s 400 4692 400 4692 0 FreeSans 600 0 0 0 A[2]
flabel metal3 s 400 3876 400 3876 0 FreeSans 600 0 0 0 A[3]
flabel metal3 s 400 3060 400 3060 0 FreeSans 600 0 0 0 A[4]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 A[5]
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 A[6]
port 7 nsew
flabel metal3 s 0 552 800 672 0 FreeSans 600 0 0 0 A[7]
port 8 nsew
flabel metal3 s 0 12792 800 12912 0 FreeSans 600 0 0 0 B[0]
port 9 nsew
flabel metal3 s 0 11976 800 12096 0 FreeSans 600 0 0 0 B[1]
port 10 nsew
flabel metal3 s 400 11220 400 11220 0 FreeSans 600 0 0 0 B[2]
flabel metal3 s 400 10404 400 10404 0 FreeSans 600 0 0 0 B[3]
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 B[4]
port 13 nsew
flabel metal3 s 400 8772 400 8772 0 FreeSans 600 0 0 0 B[5]
flabel metal3 s 0 7896 800 8016 0 FreeSans 600 0 0 0 B[6]
port 15 nsew
flabel metal3 s 400 7140 400 7140 0 FreeSans 600 0 0 0 B[7]
flabel metal5 s 1056 12672 10904 12992 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1056 9816 10904 10136 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1056 6960 10904 7280 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1056 4104 10904 4424 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal4 s 10137 2128 10457 13648 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 7699 2128 8019 13648 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 5261 2128 5581 13648 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 2823 2128 3143 13648 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal5 s 1056 12012 10904 12332 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1056 9156 10904 9476 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1056 6300 10904 6620 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1056 3444 10904 3764 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal4 s 9477 2128 9797 13648 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 7039 2128 7359 13648 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 4601 2128 4921 13648 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 2163 2128 2483 13648 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal3 s 0 15240 800 15360 0 FreeSans 600 0 0 0 opcode[0]
port 19 nsew
flabel metal3 s 0 14424 800 14544 0 FreeSans 600 0 0 0 opcode[1]
port 20 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 opcode[2]
port 21 nsew
flabel metal3 s 11200 14424 12000 14544 0 FreeSans 600 0 0 0 out[0]
port 22 nsew
flabel metal3 s 11200 12520 12000 12640 0 FreeSans 600 0 0 0 out[1]
port 23 nsew
flabel metal3 s 11200 10616 12000 10736 0 FreeSans 600 0 0 0 out[2]
port 24 nsew
flabel metal3 s 11200 8712 12000 8832 0 FreeSans 600 0 0 0 out[3]
port 25 nsew
flabel metal3 s 11200 6808 12000 6928 0 FreeSans 600 0 0 0 out[4]
port 26 nsew
flabel metal3 s 11200 4904 12000 5024 0 FreeSans 600 0 0 0 out[5]
port 27 nsew
flabel metal3 s 11200 3000 12000 3120 0 FreeSans 600 0 0 0 out[6]
port 28 nsew
flabel metal3 s 11200 1096 12000 1216 0 FreeSans 600 0 0 0 out[7]
port 29 nsew
<< properties >>
string FIXED_BBOX 0 0 12000 16000
<< end >>
