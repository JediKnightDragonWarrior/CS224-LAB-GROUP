VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lab2
  CLASS BLOCK ;
  FOREIGN lab2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 80.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END A[7]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END B[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.115 10.640 15.715 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.305 10.640 27.905 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.495 10.640 40.095 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.685 10.640 52.285 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.520 54.520 22.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 34.800 54.520 36.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.080 54.520 50.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 63.360 54.520 64.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.220 54.520 18.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 31.500 54.520 33.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.780 54.520 47.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 60.060 54.520 61.660 ;
    END
  END VPWR
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END opcode[2]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 72.120 60.000 72.720 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 62.600 60.000 63.200 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 53.080 60.000 53.680 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 43.560 60.000 44.160 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 34.040 60.000 34.640 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 24.520 60.000 25.120 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 15.000 60.000 15.600 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 5.480 60.000 6.080 ;
    END
  END out[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 54.470 68.190 ;
      LAYER li1 ;
        RECT 5.520 10.795 54.280 68.085 ;
      LAYER met1 ;
        RECT 4.210 10.640 54.670 68.240 ;
      LAYER met2 ;
        RECT 4.230 2.875 54.650 76.685 ;
      LAYER met3 ;
        RECT 4.400 75.800 56.000 76.665 ;
        RECT 3.990 73.120 56.000 75.800 ;
        RECT 4.400 71.720 55.600 73.120 ;
        RECT 3.990 69.040 56.000 71.720 ;
        RECT 4.400 67.640 56.000 69.040 ;
        RECT 3.990 64.960 56.000 67.640 ;
        RECT 4.400 63.600 56.000 64.960 ;
        RECT 4.400 63.560 55.600 63.600 ;
        RECT 3.990 62.200 55.600 63.560 ;
        RECT 3.990 60.880 56.000 62.200 ;
        RECT 4.400 59.480 56.000 60.880 ;
        RECT 3.990 56.800 56.000 59.480 ;
        RECT 4.400 55.400 56.000 56.800 ;
        RECT 3.990 54.080 56.000 55.400 ;
        RECT 3.990 52.720 55.600 54.080 ;
        RECT 4.400 52.680 55.600 52.720 ;
        RECT 4.400 51.320 56.000 52.680 ;
        RECT 3.990 48.640 56.000 51.320 ;
        RECT 4.400 47.240 56.000 48.640 ;
        RECT 3.990 44.560 56.000 47.240 ;
        RECT 4.400 43.160 55.600 44.560 ;
        RECT 3.990 40.480 56.000 43.160 ;
        RECT 4.400 39.080 56.000 40.480 ;
        RECT 3.990 36.400 56.000 39.080 ;
        RECT 4.400 35.040 56.000 36.400 ;
        RECT 4.400 35.000 55.600 35.040 ;
        RECT 3.990 33.640 55.600 35.000 ;
        RECT 3.990 32.320 56.000 33.640 ;
        RECT 4.400 30.920 56.000 32.320 ;
        RECT 3.990 28.240 56.000 30.920 ;
        RECT 4.400 26.840 56.000 28.240 ;
        RECT 3.990 25.520 56.000 26.840 ;
        RECT 3.990 24.160 55.600 25.520 ;
        RECT 4.400 24.120 55.600 24.160 ;
        RECT 4.400 22.760 56.000 24.120 ;
        RECT 3.990 20.080 56.000 22.760 ;
        RECT 4.400 18.680 56.000 20.080 ;
        RECT 3.990 16.000 56.000 18.680 ;
        RECT 4.400 14.600 55.600 16.000 ;
        RECT 3.990 11.920 56.000 14.600 ;
        RECT 4.400 10.520 56.000 11.920 ;
        RECT 3.990 7.840 56.000 10.520 ;
        RECT 4.400 6.480 56.000 7.840 ;
        RECT 4.400 6.440 55.600 6.480 ;
        RECT 3.990 5.080 55.600 6.440 ;
        RECT 3.990 3.760 56.000 5.080 ;
        RECT 4.400 2.895 56.000 3.760 ;
  END
END lab2
END LIBRARY

